0.507218	0.494949	0.486663	0.308828
0.500678	0.587537	0.664670	0.429262
0.527465	0.598560	0.527895	0.295296
0.527966	0.388086	0.410960	0.354974
0.544203	0.428920	0.599219	0.345108
0.564248	0.385916	0.370601	0.385039
0.560935	0.575417	0.415849	0.376575
0.577571	0.597395	0.408281	0.473651
0.576304	0.498664	0.360713	0.371034
0.546683	0.545423	0.473409	0.452635
0.632409	0.625542	0.587933	0.367366
0.570873	0.425262	0.632359	0.493018
0.569296	0.504110	0.496267	0.350804
0.571996	0.505503	0.514490	0.341455
0.504371	0.593184	0.474356	0.289583
0.509895	0.469301	0.312361	0.347802
0.588081	0.520679	0.451081	0.400045
0.574765	0.574970	0.402260	0.386736
0.502227	0.469874	0.533935	0.366580
0.524331	0.453641	0.405218	0.330668
0.517153	0.440760	0.457895	0.372519
0.530644	0.510915	0.393348	0.417545
0.584106	0.559858	0.578996	0.342832
0.552836	0.555891	0.481003	0.384248
0.562160	0.476098	0.443729	0.399493
0.600889	0.539802	0.263843	0.456541
0.530923	0.460615	0.419672	0.395465
0.561792	0.555444	0.525129	0.438325
0.577032	0.504151	0.408098	0.367119
0.495427	0.556791	0.484364	0.310131
0.523320	0.463306	0.410345	0.480305
0.565056	0.460128	0.494211	0.475645
0.606674	0.564577	0.274779	0.450504
0.580113	0.463369	0.366760	0.407662
0.536838	0.418381	0.441862	0.405584
0.554402	0.606853	0.621059	0.389695
0.621639	0.464961	0.435688	0.408811
0.572213	0.435921	0.540103	0.406130
0.553856	0.477450	0.490768	0.415067
0.526873	0.539897	0.383454	0.353629
0.565219	0.514931	0.491413	0.351506
0.467107	0.561382	0.443587	0.308652
0.492949	0.525333	0.510924	0.347194
0.588560	0.539582	0.765336	0.389430
0.492792	0.421744	0.308385	0.305626
0.577378	0.592894	0.428020	0.372156
0.591103	0.441996	0.487685	0.448798
0.563393	0.452565	0.249209	0.409664
0.508324	0.549465	0.272427	0.416632
0.583214	0.443639	0.405305	0.387962
0.542423	0.446758	0.321762	0.378280
0.730681	0.513707	0.434146	0.451108
0.594459	0.450380	0.311672	0.452428
0.597823	0.457650	0.400483	0.393513
0.557161	0.463081	0.471805	0.357191
0.542091	0.443834	0.540603	0.397069
0.542837	0.499593	0.163108	0.333269
0.529535	0.524810	0.218462	0.407939
0.622537	0.501100	0.741571	0.412018
0.535382	0.463487	0.494433	0.465035
0.493629	0.522116	0.406437	0.327724
0.590530	0.496306	0.205456	0.362333
0.572438	0.451610	0.446586	0.359574
0.600755	0.491348	0.282712	0.393860
0.524836	0.476953	0.497962	0.398321
0.508585	0.422206	0.506470	0.350777
0.571426	0.583605	0.234386	0.518727
0.588841	0.489005	0.205901	0.372552
0.546730	0.642539	0.403710	0.353405
0.568952	0.469532	0.425421	0.423356
0.600953	0.476186	0.398611	0.473420
0.593394	0.638757	0.508924	0.394751
0.581779	0.653903	0.494697	0.324451
0.584121	0.522436	0.571998	0.357613
0.509417	0.506136	0.402132	0.426233
0.631997	0.438358	0.502832	0.405494
0.465870	0.584118	0.451386	0.268141
0.527922	0.390285	0.395139	0.384743
0.556421	0.475088	0.640916	0.360214
0.561673	0.534732	0.418789	0.382538
0.579903	0.548831	0.582476	0.350420
0.620847	0.637031	0.600750	0.428535
0.663089	0.422814	0.442116	0.425304
0.591339	0.571016	0.308775	0.334922
0.492084	0.485067	0.384248	0.428355
0.545677	0.452074	0.428627	0.428418
0.597916	0.434950	0.440570	0.461763
0.469430	0.488470	0.398758	0.295887
0.528447	0.587804	0.789025	0.353410
0.541678	0.501669	0.598813	0.370948
0.489907	0.517767	0.502323	0.331069
0.573975	0.623398	0.523294	0.352725
0.546526	0.401637	0.291932	0.364181
0.551143	0.565267	0.544477	0.383874
0.636052	0.398080	0.484273	0.406751
0.583457	0.601944	0.542017	0.411397
0.667924	0.555115	0.518213	0.407316
0.556503	0.436633	0.322443	0.373714
0.545042	0.481994	0.459324	0.355459
0.548033	0.540306	0.605424	0.389053
0.562487	0.593475	0.391613	0.468597
0.597827	0.483310	0.374478	0.481505
0.540252	0.440664	0.457199	0.365489
0.574173	0.449763	0.642490	0.383828
0.579596	0.537192	0.287393	0.442235
0.528789	0.569535	0.552774	0.368344
0.569201	0.454860	0.324792	0.406626
0.560940	0.604588	0.575837	0.357356
0.515537	0.520308	0.483984	0.452068
0.504210	0.445975	0.598937	0.414684
0.536217	0.510896	0.507854	0.416450
0.585426	0.534425	0.535479	0.442669
0.553701	0.439972	0.695700	0.365509
0.589733	0.597807	0.495533	0.363295
0.534393	0.431851	0.341018	0.339046
0.617798	0.506887	0.529353	0.449171
0.524620	0.609270	0.307778	0.365247
0.591435	0.500680	0.416008	0.415711
0.577879	0.440439	0.569942	0.411466
0.516297	0.573096	0.280873	0.300782
0.471969	0.595976	0.497108	0.473889
0.547009	0.467059	0.144963	0.368014
0.620188	0.506427	0.391398	0.471387
0.566094	0.575626	0.551269	0.336565
0.548357	0.552442	0.433769	0.364930
0.531322	0.532799	0.873106	0.315591
0.624875	0.455966	0.422429	0.501826
0.627398	0.475870	0.547490	0.467218
0.522477	0.599816	0.409924	0.296929
0.522829	0.433813	0.335401	0.388581
0.535832	0.391745	0.341883	0.337017
0.582700	0.549921	0.345823	0.430812
0.586475	0.568193	0.677598	0.343752
0.493442	0.577222	0.267857	0.419648
0.590571	0.542303	0.697339	0.517327
0.536247	0.492944	0.452467	0.417559
0.504568	0.566903	0.343938	0.331497
0.476114	0.540893	0.484502	0.302122
0.564987	0.573903	0.407345	0.467108
0.546097	0.495385	0.564890	0.373061
0.563033	0.525019	0.588337	0.345772
0.539115	0.498123	0.400543	0.336759
0.588908	0.543673	0.462060	0.391812
0.581948	0.421727	0.588192	0.470192
0.597121	0.479895	0.411266	0.409867
0.594670	0.620614	0.724509	0.465073
0.528120	0.412911	0.673638	0.409194
0.588637	0.463714	0.297525	0.407594
0.583956	0.534789	0.390189	0.352037
0.583847	0.525518	0.794414	0.632157
0.634483	0.494032	0.527442	0.454300
0.544429	0.530073	0.317801	0.349156
0.561171	0.537040	0.644220	0.503480
0.547395	0.533091	0.521455	0.379043
0.516277	0.651606	0.320559	0.479041
0.592782	0.521912	0.470610	0.391287
0.566103	0.521714	0.701508	0.358344
0.569478	0.586859	0.484287	0.397510
0.509770	0.515909	0.653549	0.461021
0.529977	0.555454	0.429977	0.319503
0.557945	0.410170	0.329208	0.369770
0.459936	0.456636	0.264521	0.375620
0.464681	0.610956	0.589108	0.293525
0.568548	0.542676	0.359013	0.362296
0.512079	0.495930	0.299109	0.359183
0.636469	0.461132	0.369891	0.501359
0.506659	0.478183	0.511575	0.482927
0.588558	0.465044	0.322337	0.351270
0.524633	0.481174	0.603630	0.318201
0.671638	0.537146	0.372743	0.420149
0.634922	0.614105	0.377526	0.525522
0.535525	0.447422	0.367612	0.390006
0.580277	0.591500	0.537464	0.341106
0.506751	0.517151	0.320032	0.467596
0.503099	0.443191	0.362904	0.406602
0.606949	0.551956	0.647366	0.435090
0.568510	0.444224	0.489795	0.422180
0.551439	0.467843	0.306453	0.403762
0.535340	0.501918	0.291224	0.342231
0.640805	0.481188	0.475832	0.394197
0.497311	0.512749	0.542918	0.341402
0.527415	0.427747	0.405596	0.449183
0.544131	0.468800	0.709503	0.333794
0.584196	0.548511	0.573423	0.345014
0.538218	0.612485	0.555461	0.333982
0.536867	0.551190	0.489059	0.391164
0.598848	0.367603	0.464116	0.395247
0.590764	0.474661	0.637389	0.395340
0.646118	0.506508	0.621459	0.459643
0.570079	0.480529	0.428380	0.344265
0.610459	0.438533	0.686542	0.379604
0.615357	0.411629	0.252755	0.390695
0.583188	0.470364	0.410463	0.422414
0.567054	0.516298	0.448553	0.358916
0.448077	0.574960	0.509685	0.268698
0.559923	0.688850	0.516771	0.459060
0.525652	0.609665	0.284701	0.349840
0.679543	0.549426	0.564320	0.399269
0.647689	0.629511	0.417244	0.467482
0.590828	0.475393	0.376707	0.490259
0.493346	0.458359	0.589833	0.395799
0.563939	0.403408	0.381282	0.508312
0.592826	0.577683	0.194398	0.412079
0.571955	0.415657	0.414466	0.400291
0.550814	0.591077	0.389287	0.485089
0.486712	0.427623	0.411068	0.424002
0.525473	0.515797	0.509156	0.360663
0.557497	0.452674	0.437008	0.475262
0.535328	0.361854	0.342875	0.458926
0.571369	0.478719	0.736774	0.372322
0.509516	0.467927	0.246051	0.333865
0.541914	0.592516	0.345335	0.311224
0.602917	0.481728	0.874596	0.433279
0.475498	0.431476	0.443784	0.353639
0.621257	0.550996	0.599823	0.469671
0.537873	0.497590	0.517155	0.383156
0.480366	0.546579	0.428577	0.320865
0.599177	0.461098	0.372945	0.363569
0.571104	0.458467	0.370095	0.416615
0.664373	0.501965	0.576110	0.441249
0.498694	0.470485	0.723733	0.342085
0.608652	0.341178	0.572678	0.459828
0.606375	0.606990	0.562828	0.345225
0.535505	0.457915	0.408661	0.331020
0.519104	0.565699	0.352981	0.335869
0.553092	0.478025	0.500684	0.364128
0.582785	0.568210	0.661686	0.342889
0.498619	0.542789	0.519009	0.289117
0.601056	0.547911	0.452695	0.356179
0.500182	0.579221	0.453288	0.465042
0.610101	0.653653	0.621037	0.354000
0.593264	0.334818	0.414771	0.382157
0.537967	0.569044	0.734339	0.376873
0.587200	0.547352	0.553298	0.358283
0.561408	0.497292	0.718482	0.355767
0.508963	0.542763	0.610018	0.408147
0.545676	0.573941	0.586553	0.325263
0.474129	0.588374	0.302102	0.289646
0.565712	0.513130	0.606073	0.411090
0.603563	0.491795	0.416165	0.419505
0.623580	0.573396	0.322086	0.429024
0.607406	0.639838	0.315037	0.350708
0.670953	0.535164	0.226855	0.438694
0.577650	0.462275	0.510745	0.367709
0.586943	0.517999	0.300665	0.363901
0.551712	0.526698	0.494060	0.327796
0.487813	0.450546	0.432324	0.416668
0.594636	0.611708	0.485741	0.393789
0.607269	0.607883	0.533074	0.383884
0.527763	0.464911	0.592375	0.452829
0.553247	0.364024	0.428618	0.362224
0.510576	0.569251	0.595206	0.330735
0.563061	0.372506	0.398140	0.355138
0.605817	0.454517	0.620279	0.366254
0.540228	0.529115	0.519904	0.514848
0.491920	0.501049	0.506103	0.340863
0.529476	0.472320	0.530978	0.352875
0.543737	0.566883	0.393202	0.370153
0.568258	0.634940	0.092661	0.352562
0.525549	0.467872	0.535166	0.379252
0.525501	0.474799	0.499952	0.417331
0.540669	0.434134	0.590371	0.369689
0.599289	0.459085	0.183154	0.404587
0.409121	0.616328	0.292255	0.375557
0.573146	0.469828	0.287703	0.376725
0.552168	0.542883	0.530115	0.380746
0.621320	0.534888	0.721567	0.465447
0.580112	0.522750	0.518452	0.405438
0.542601	0.393904	0.428917	0.386766
0.525195	0.525380	0.225866	0.342502
0.532286	0.551935	0.357335	0.376760
0.557919	0.557305	0.497518	0.414071
0.509427	0.471543	0.387616	0.444154
0.602968	0.482520	0.106127	0.373115
0.549912	0.535403	0.375494	0.370284
0.574565	0.535693	0.430694	0.359078
0.576145	0.573450	0.334846	0.414907
0.496671	0.572221	0.373856	0.349347
0.558942	0.506309	0.788310	0.425705
0.556677	0.478984	0.742991	0.412802
0.567156	0.420943	0.558534	0.365887
0.512911	0.514672	0.378099	0.402347
0.540728	0.622866	0.430073	0.366739
0.552180	0.509805	0.437275	0.371867
0.577450	0.498112	0.178854	0.414514
0.579706	0.534846	0.213286	0.390349
0.575176	0.473135	0.362757	0.401730
0.510076	0.483268	0.381540	0.359672
0.580830	0.436919	0.277438	0.403029
0.550071	0.616397	0.514303	0.446846
0.609174	0.357168	0.340523	0.386327
0.573471	0.538338	0.436314	0.362425
0.556413	0.451612	0.351444	0.368663
0.619673	0.476522	0.404022	0.372479
0.616165	0.648148	0.491367	0.378276
0.522250	0.531701	0.409766	0.479801
0.539310	0.517053	0.495082	0.321205
0.506388	0.422008	0.288729	0.342820
0.530734	0.581397	0.085859	0.346699
0.514894	0.462008	0.530938	0.420710
0.490249	0.652116	0.193443	0.342137
0.535252	0.522138	0.683340	0.446629
0.591339	0.533714	0.371654	0.392920
0.563671	0.593005	0.523869	0.390099
0.543071	0.498092	0.454343	0.345588
0.498138	0.615087	0.587563	0.396873
0.539699	0.477604	0.521222	0.395530
0.534000	0.481148	0.367115	0.354371
0.501515	0.519018	0.707288	0.492027
0.570402	0.503645	0.616461	0.384864
0.575836	0.398556	0.634914	0.420171
0.628730	0.539224	0.333885	0.402471
0.511032	0.635721	0.342215	0.335719
0.505985	0.641879	0.531658	0.343125
0.559720	0.524967	0.432212	0.374445
0.512890	0.420743	0.399027	0.419920
0.566901	0.522110	0.380303	0.434078
0.514475	0.496283	0.124016	0.478591
0.586917	0.502295	0.589985	0.362396
0.542282	0.536607	0.172261	0.345634
0.619684	0.610538	0.582021	0.440328
0.478095	0.530905	0.667079	0.300844
0.554142	0.518672	0.256552	0.426093
0.516400	0.524416	0.564944	0.440835
0.670532	0.418241	0.502726	0.499757
0.519327	0.653993	0.257392	0.325468
0.578181	0.479055	0.636703	0.347244
0.604846	0.562739	0.230065	0.365330
0.526982	0.544972	0.531854	0.323600
0.555018	0.710519	0.680832	0.410787
0.525152	0.497190	0.309269	0.307218
0.530325	0.472157	0.488978	0.455570
0.606121	0.550982	0.529182	0.358090
0.526187	0.566755	0.410705	0.377964
0.579157	0.536841	0.468034	0.445635
0.558548	0.451738	0.528954	0.450843
0.568424	0.485638	0.588866	0.498633
0.609395	0.437063	0.549729	0.512237
0.620429	0.440143	0.345882	0.453458
0.475109	0.543022	0.368591	0.369191
0.488990	0.548154	0.410484	0.305380
0.466839	0.510968	0.617703	0.327029
0.487635	0.484145	0.445472	0.374994
0.561661	0.500751	0.532081	0.383925
0.563140	0.498308	0.407372	0.382228
0.506732	0.577660	0.383982	0.354283
0.551277	0.637136	0.604175	0.503678
0.575038	0.464744	0.295559	0.357509
0.549891	0.396971	0.640655	0.360232
0.524735	0.553276	0.322978	0.303160
0.527385	0.338814	0.459003	0.420848
0.537192	0.452672	0.548660	0.354616
0.526288	0.463430	0.742066	0.337072
0.568814	0.492480	0.322880	0.371042
0.603756	0.524747	0.462038	0.446231
0.570023	0.537264	0.656539	0.364034
0.539926	0.449374	0.480748	0.405955
0.534421	0.450319	0.458204	0.377115
0.540056	0.546864	0.409492	0.416338
0.571034	0.414439	0.326214	0.494176
0.543536	0.632152	0.513559	0.378089
0.545769	0.386921	0.471977	0.348222
0.595356	0.413962	0.437389	0.407611
0.614448	0.509001	0.798454	0.400366
0.597537	0.589994	0.517414	0.367196
0.561378	0.590456	0.680398	0.483665
0.611382	0.554362	0.114282	0.426524
0.547326	0.489822	0.299964	0.349723
0.524830	0.479739	0.472907	0.418579
0.607939	0.544037	0.245984	0.366387
0.576640	0.553997	0.428482	0.375616
0.554991	0.512301	0.626981	0.349561
0.537944	0.568680	0.153487	0.457325
0.551877	0.494193	0.371891	0.326633
0.531087	0.470330	0.291593	0.387649
0.580960	0.551489	0.433195	0.393349
0.546491	0.433859	0.784952	0.458418
0.592436	0.552519	0.562308	0.417260
0.605669	0.428255	0.188423	0.368278
0.474380	0.564546	0.557114	0.368639
0.607337	0.566242	0.756810	0.415908
0.515666	0.518747	0.499739	0.375505
0.551531	0.358283	0.538768	0.514424
0.552911	0.543204	0.431343	0.389644
0.542011	0.509453	0.287408	0.362796
0.571980	0.431113	0.425372	0.472802
0.505349	0.528502	0.285498	0.345019
0.489855	0.477309	0.382206	0.384917
0.549905	0.396559	0.579581	0.423488
0.578394	0.418878	0.151246	0.388564
0.658724	0.441271	0.204459	0.417646
0.563170	0.474115	0.210469	0.413993
0.596530	0.473630	0.271688	0.390266
0.581325	0.537105	0.391646	0.431766
0.578662	0.484999	0.627870	0.345723
0.540192	0.497607	0.286534	0.361175
0.585388	0.503414	0.630843	0.402458
0.605245	0.457596	0.350639	0.407729
0.537865	0.539748	0.434625	0.313081
0.626669	0.531046	0.540986	0.501494
0.619647	0.586618	0.232853	0.390634
0.649173	0.601721	0.620147	0.370462
0.574355	0.552998	0.636755	0.372378
0.554295	0.398644	0.232276	0.385875
0.536862	0.431631	0.409309	0.475112
0.546038	0.500870	0.599304	0.404369
0.634747	0.562411	0.557798	0.364894
0.603810	0.525336	0.646069	0.362485
0.655360	0.483695	0.389741	0.438923
0.612264	0.562547	0.352325	0.444877
0.530645	0.497306	0.324986	0.394461
0.577061	0.426127	0.354371	0.414248
0.567296	0.539821	0.363203	0.357868
0.553500	0.459041	0.384776	0.349996
0.583184	0.606792	0.569614	0.342100
0.594584	0.544415	0.392217	0.426759
0.581474	0.476023	0.483080	0.398555
0.559026	0.656776	0.276586	0.407888
0.503839	0.604087	0.545557	0.333308
0.504592	0.566992	0.682051	0.320719
0.551846	0.393131	0.359621	0.367196
0.630139	0.601054	0.404787	0.457805
0.618800	0.330848	0.557198	0.439701
0.643152	0.546240	0.219583	0.376892
0.519417	0.539030	0.283398	0.357867
0.544181	0.672040	0.227899	0.361744
0.663015	0.449696	0.393183	0.483844
0.568623	0.505477	0.341343	0.335316
0.585218	0.548826	0.492956	0.345595
0.607124	0.609182	0.546352	0.342313
0.592257	0.351957	0.629298	0.541281
0.504760	0.549026	0.256551	0.464740
0.576135	0.606094	0.352561	0.374070
0.538179	0.561873	0.402285	0.359391
0.571565	0.531765	0.528707	0.334594
0.570349	0.465078	0.554425	0.416760
0.588742	0.555078	0.440598	0.343252
0.541808	0.405239	0.354865	0.391510
0.528731	0.526219	0.394363	0.322712
0.537033	0.624137	0.345286	0.366432
0.539101	0.519849	0.411290	0.350230
0.488838	0.482352	0.296757	0.403348
0.568882	0.496643	0.392179	0.339493
0.609854	0.624353	0.301703	0.393850
0.589822	0.501907	0.659036	0.386074
0.523727	0.466964	0.341361	0.403216
0.544930	0.520823	0.695659	0.333209
0.531828	0.464726	0.264854	0.321570
0.539706	0.444255	0.569199	0.371687
0.502150	0.535495	0.392867	0.416838
0.547434	0.628552	0.659961	0.318173
0.604312	0.421620	0.461602	0.382682
0.540641	0.439101	0.575174	0.407156
0.505762	0.268167	0.399911	0.455632
0.576159	0.480474	0.384070	0.389192
0.546529	0.628329	0.494162	0.461872
0.560339	0.503678	0.567856	0.388419
0.572841	0.482717	0.514150	0.398830
0.528807	0.535216	0.594608	0.323896
0.455187	0.601436	0.371603	0.354181
0.481886	0.488823	0.640349	0.398048
0.605979	0.408516	0.265944	0.399958
0.588896	0.455780	0.520143	0.447349
0.485970	0.550219	0.642864	0.484740
0.541808	0.554823	0.317968	0.493654
0.538922	0.529307	0.534958	0.476532
0.656180	0.531444	0.426188	0.460852
0.550135	0.588263	0.338529	0.410133
0.539058	0.514909	0.224518	0.385846
0.593730	0.522844	0.615529	0.353871
0.641091	0.683437	0.487174	0.351760
0.572300	0.430206	0.308532	0.355717
0.598332	0.456610	0.475942	0.399684
0.548432	0.569654	0.435318	0.440385
0.646901	0.511394	0.463098	0.423622
0.611794	0.518767	0.396965	0.442291
0.529499	0.415780	0.652876	0.331192
0.543856	0.371660	0.252466	0.431340
0.589422	0.499083	0.651244	0.384539
0.473382	0.392049	0.341011	0.472458
0.565520	0.497839	0.388301	0.375439
0.529933	0.563411	0.293658	0.407364
0.598997	0.403200	0.326335	0.427086
0.580759	0.483751	0.577802	0.386713
0.495018	0.518538	0.451151	0.328902
0.519670	0.543127	0.316441	0.392064
0.589950	0.482878	0.685896	0.418447
0.597863	0.522752	0.458482	0.427461
0.610811	0.449603	0.531900	0.385374
0.640771	0.460626	0.247879	0.445394
0.527353	0.570539	0.422389	0.397805
0.561995	0.579035	0.368180	0.371266
0.571749	0.682489	0.442915	0.343258
0.577138	0.509015	0.410700	0.464163
0.621146	0.433271	0.350896	0.383459
0.488054	0.450223	0.387976	0.389770
0.554458	0.569349	0.605631	0.479099
0.544266	0.572662	0.255554	0.427542
0.578963	0.522533	0.446522	0.502981
0.536429	0.531890	0.612074	0.335199
0.608750	0.524743	0.430057	0.378767
0.614996	0.430251	0.431945	0.428250
0.580067	0.653570	0.415523	0.323936
0.489805	0.583126	0.346109	0.327556
0.590595	0.362541	0.584915	0.389777
0.514908	0.449308	0.191814	0.357490
0.550405	0.538628	0.528292	0.338229
0.477574	0.470989	0.450032	0.386468
0.593698	0.607928	0.330306	0.417786
0.564318	0.428303	0.486222	0.348257
0.545434	0.494988	0.470916	0.375125
0.572820	0.500644	0.535756	0.359176
0.579919	0.544242	0.360610	0.346400
0.514749	0.591615	0.434742	0.334466
0.534924	0.412216	0.480096	0.423614
0.504770	0.460835	0.437620	0.356907
0.602252	0.425302	0.431938	0.404198
0.479374	0.626555	0.558267	0.298910
0.554808	0.666010	0.402078	0.383853
0.593948	0.550938	0.471237	0.350769
0.543202	0.545003	0.273274	0.432580
0.633867	0.498909	0.327928	0.395733
0.532476	0.464567	0.269304	0.415562
0.503772	0.549988	0.280824	0.457651
0.500475	0.503994	0.428790	0.376996
0.580306	0.479032	0.445482	0.445931
0.481589	0.593893	0.749835	0.456110
0.613677	0.457547	0.520556	0.488406
0.588833	0.514777	0.276578	0.423788
0.538113	0.500062	0.416029	0.338303
0.482119	0.476012	0.713341	0.343541
0.535029	0.592781	0.427016	0.310947
0.615488	0.521682	0.700471	0.372542
0.504706	0.519657	0.636364	0.412670
0.490002	0.443343	0.418882	0.472665
0.514363	0.635205	0.240881	0.355908
0.564785	0.567556	0.454000	0.517513
0.580307	0.617298	0.446365	0.452674
0.522872	0.679577	0.496640	0.326444
0.520490	0.535841	0.541744	0.325849
0.546100	0.508507	0.586993	0.326516
0.602889	0.329551	0.583996	0.428301
0.556767	0.464918	0.639641	0.466650
0.553673	0.527063	0.299016	0.390238
0.582291	0.547286	0.310271	0.591673
0.629164	0.443130	0.370383	0.409460
0.625776	0.556311	0.500024	0.385410
0.551203	0.368272	0.701300	0.465925
0.556415	0.634811	0.744057	0.335908
0.613506	0.560273	0.640873	0.374826
0.554857	0.480761	0.508844	0.406142
0.616373	0.526968	0.449750	0.418721
0.597188	0.501246	0.609519	0.467396
0.507357	0.498423	0.393670	0.305201
0.599792	0.504264	0.462313	0.408655
0.600118	0.436098	0.686233	0.370311
0.592043	0.517997	0.469606	0.403131
0.522827	0.492263	0.396188	0.367906
0.598424	0.570974	0.470287	0.441945
0.521958	0.450476	0.416470	0.399870
0.568412	0.573173	0.486069	0.415976
0.556788	0.552465	0.403072	0.407748
0.573775	0.450842	0.314289	0.460535
0.656477	0.740957	0.196097	0.391068
0.571823	0.448034	0.358887	0.360638
0.590240	0.576359	0.439729	0.504971
0.634569	0.519423	0.306516	0.435171
0.529122	0.483978	0.397355	0.343073
0.630960	0.545332	0.405087	0.380823
0.605043	0.501703	0.425440	0.428172
0.489091	0.472089	0.294214	0.325635
0.572803	0.423623	0.497869	0.359985
0.600414	0.496424	0.213662	0.416682
0.477794	0.444829	0.362241	0.473775
0.617696	0.453092	0.650340	0.376123
0.536109	0.418156	0.538290	0.363804
0.599860	0.467723	0.442429	0.449242
0.589169	0.562001	0.277423	0.365049
0.526729	0.528087	0.400301	0.441234
0.535316	0.412879	0.599975	0.332123
0.552036	0.591181	0.579709	0.327342
0.576742	0.520181	0.504558	0.394229
0.543597	0.483647	0.384157	0.354267
0.547190	0.501775	0.457747	0.368134
0.501317	0.584009	0.678056	0.317552
0.458631	0.364252	0.533097	0.312061
0.550826	0.582597	0.277877	0.321477
0.582683	0.524750	0.325563	0.351248
0.560262	0.482915	0.409435	0.485883
0.519671	0.635177	0.640435	0.343702
0.603348	0.425515	0.360886	0.382152
0.576228	0.417011	0.444196	0.401275
0.533481	0.420425	0.255025	0.325742
0.568667	0.493639	0.301273	0.351914
0.571551	0.497741	0.576107	0.598342
0.475825	0.395512	0.261509	0.386070
0.529671	0.398472	0.454794	0.357475
0.513851	0.542242	0.535023	0.373090
0.538975	0.536615	0.474869	0.343535
0.636572	0.557952	0.431131	0.402022
0.593604	0.511875	0.427111	0.448364
0.540801	0.412569	0.449193	0.372023
0.585773	0.501221	0.473135	0.391216
0.559349	0.526863	0.147858	0.346104
0.525733	0.376208	0.550776	0.351439
0.609961	0.302504	0.528302	0.400252
0.582658	0.553062	0.395076	0.421076
0.491950	0.618216	0.522054	0.408592
0.630562	0.629319	0.468610	0.426748
0.615709	0.458995	0.458141	0.448940
0.587052	0.346313	0.428088	0.413659
0.605033	0.644681	0.523589	0.352913
0.604398	0.667275	0.501540	0.465307
0.593490	0.527094	0.375667	0.366534
0.572101	0.656925	0.333929	0.537571
0.635912	0.430224	0.364945	0.444545
0.648603	0.594079	0.574212	0.404544
0.516368	0.567465	0.462567	0.434269
0.560947	0.330321	0.476645	0.361525
0.576131	0.495816	0.524056	0.411880
0.531188	0.361362	0.262234	0.362424
0.514728	0.478189	0.272509	0.321869
0.541921	0.613345	0.440484	0.394628
0.604389	0.619427	0.622881	0.342698
0.517389	0.432014	0.445244	0.368156
0.583301	0.423960	0.250764	0.471301
0.548945	0.462470	0.257243	0.381141
0.547301	0.432472	0.472948	0.480610
0.557532	0.449312	0.442144	0.481972
0.599748	0.511832	0.243317	0.402212
0.539593	0.506813	0.528867	0.360658
0.515592	0.541085	0.455669	0.331098
0.626442	0.652539	0.358992	0.374164
0.601798	0.535279	0.635305	0.418336
0.614069	0.457079	0.228416	0.369251
0.599031	0.543035	0.587209	0.464222
0.640737	0.588467	0.508331	0.426864
0.546476	0.585931	0.548976	0.320957
0.556067	0.487786	0.522959	0.344141
0.606285	0.414035	0.131172	0.455439
0.611243	0.618315	0.477170	0.355415
0.567622	0.529692	0.423904	0.404778
0.523467	0.423001	0.320852	0.369297
0.460144	0.445551	0.455084	0.346255
0.568865	0.632789	0.503888	0.396532
0.549232	0.516609	0.713934	0.324297
0.524890	0.556095	0.501485	0.367685
0.584168	0.392740	0.315136	0.444489
0.599570	0.601454	0.589237	0.346195
0.518254	0.598840	0.541858	0.412968
0.591215	0.465033	0.524148	0.357168
0.498341	0.645389	0.683622	0.402264
0.585442	0.384581	0.450605	0.389471
0.626882	0.570625	0.298291	0.449032
0.550685	0.586490	0.451194	0.358621
0.577052	0.595256	0.349515	0.324990
0.536359	0.480533	0.482833	0.408610
0.546383	0.508671	0.362057	0.412241
0.574867	0.565141	0.531014	0.335706
0.480119	0.541434	0.386987	0.395474
0.530453	0.571988	0.364927	0.314115
0.578093	0.569966	0.216477	0.456038
0.552620	0.373847	0.401550	0.389981
0.579044	0.372615	0.345520	0.447123
0.572493	0.550216	0.666720	0.417527
0.623903	0.576014	0.556565	0.376232
0.615724	0.482135	0.284484	0.431794
0.519400	0.610446	0.470125	0.424854
0.509621	0.528848	0.579438	0.386518
0.654849	0.537861	0.761616	0.460502
0.531742	0.614031	0.336106	0.313072
0.549722	0.593624	0.549291	0.374810
0.516782	0.644359	0.440523	0.316245
0.575298	0.531099	0.769969	0.400310
0.453861	0.489434	0.440245	0.414154
0.556980	0.428081	0.490858	0.384154
0.502253	0.582501	0.298370	0.282855
0.633425	0.517908	0.300442	0.422709
0.589504	0.427511	0.554003	0.372089
0.538985	0.571085	0.602274	0.414430
0.537297	0.525862	0.612209	0.436720
0.556251	0.555640	0.615232	0.384838
0.611509	0.527812	0.373330	0.405901
0.558191	0.416810	0.505886	0.419803
0.560922	0.524998	0.434908	0.349478
0.557012	0.431112	0.409117	0.356335
0.572170	0.712517	0.341769	0.407590
0.586449	0.480588	0.327951	0.447609
0.572652	0.519462	0.271562	0.389481
0.522261	0.551204	0.648839	0.367546
0.526871	0.559126	0.182885	0.373380
0.527455	0.532548	0.520435	0.335992
0.581881	0.539847	0.325899	0.482990
0.581058	0.421357	0.360275	0.432132
0.514063	0.510702	0.277312	0.449713
0.563242	0.564166	0.447445	0.325650
0.454933	0.554410	0.515796	0.325347
0.576116	0.523685	0.400412	0.410672
0.526160	0.483092	0.508063	0.354092
0.555349	0.579293	0.437000	0.355692
0.557603	0.645085	0.479155	0.365409
0.570911	0.458710	0.234495	0.415302
0.661601	0.587100	0.472705	0.393372
0.507962	0.475352	0.610348	0.377287
0.514700	0.431247	0.482446	0.379874
0.528645	0.426073	0.653337	0.337458
0.593636	0.531761	0.500349	0.363970
0.595499	0.502874	0.571308	0.478039
0.583417	0.452734	0.400761	0.368852
0.631547	0.537870	0.349146	0.366025
0.569836	0.555876	0.539923	0.388629
0.629591	0.536173	0.382330	0.380987
0.612829	0.650596	0.455939	0.351925
0.582939	0.397038	0.248111	0.383457
0.590589	0.546137	0.441069	0.453542
0.570665	0.546029	0.501668	0.341874
0.492572	0.485324	0.191241	0.401369
0.564956	0.562787	0.437564	0.350919
0.560338	0.458963	0.351684	0.410148
0.560268	0.410069	0.555401	0.443494
0.531066	0.393732	0.614313	0.350375
0.537151	0.552956	0.392119	0.456960
0.565487	0.557671	0.381166	0.355266
0.484991	0.513247	0.502359	0.366718
0.558342	0.491474	0.058465	0.409502
0.556641	0.566824	0.437933	0.351711
0.583611	0.563841	0.311772	0.347394
0.609167	0.545651	0.441929	0.490504
0.603114	0.413402	0.388344	0.474598
0.546921	0.549029	0.298796	0.386729
0.547293	0.560116	0.380455	0.380812
0.563780	0.587129	0.540361	0.318208
0.545719	0.449317	0.319280	0.327302
0.599928	0.474443	0.408979	0.421819
0.459511	0.356259	0.351623	0.392954
0.557867	0.411210	0.327441	0.344558
0.502606	0.449911	0.450301	0.371666
0.503862	0.483688	0.322513	0.330115
0.646206	0.523797	0.595365	0.448913
0.545882	0.533560	0.579451	0.395015
0.583876	0.519061	0.542321	0.384857
0.588488	0.351126	0.365531	0.444723
0.586492	0.488060	0.338913	0.437378
0.612963	0.452378	0.424255	0.401460
0.631191	0.551105	0.475338	0.434842
0.653978	0.504327	0.430021	0.441374
0.550729	0.462487	0.317051	0.355927
0.545644	0.486550	0.470569	0.350755
0.493235	0.637394	0.313210	0.309393
0.588910	0.614580	0.362801	0.337592
0.549343	0.378624	0.720212	0.390102
0.574060	0.527879	0.481076	0.422363
0.631796	0.583086	0.178639	0.405808
0.579702	0.548893	0.592448	0.371977
0.560973	0.375975	0.494460	0.352939
0.502154	0.518688	0.454206	0.507377
0.533727	0.477730	0.581359	0.387106
0.566949	0.546671	0.409437	0.365349
0.563916	0.477088	0.606902	0.432777
0.542125	0.479178	0.515660	0.346154
0.585148	0.421288	0.400726	0.361053
0.582273	0.406072	0.477153	0.379851
0.520320	0.644762	0.373643	0.294779
0.508665	0.499464	0.556365	0.433830
0.621771	0.643253	0.592173	0.431009
0.533994	0.423035	0.597422	0.395582
0.573761	0.462682	0.463202	0.433979
0.553810	0.388867	0.322053	0.403988
0.481198	0.459163	0.137337	0.306137
0.492969	0.540808	0.322161	0.296810
0.529561	0.577869	0.582950	0.421375
0.494404	0.631166	0.434304	0.336645
0.497820	0.613858	0.559797	0.305985
0.586879	0.692026	0.440948	0.351668
0.669884	0.478414	0.431722	0.463517
0.492886	0.501730	0.440603	0.440222
0.556629	0.559319	0.364620	0.400308
0.519506	0.365670	0.292305	0.327378
0.538129	0.556376	0.491760	0.308922
0.561285	0.373222	0.264730	0.374282
0.540711	0.551221	0.544149	0.351620
0.500391	0.587521	0.387974	0.363652
0.627954	0.614793	0.385967	0.362924
0.546383	0.455977	0.368461	0.373980
0.525541	0.584957	0.485834	0.409024
0.573891	0.488628	0.461915	0.477909
0.666331	0.409089	0.578786	0.472998
0.590963	0.489321	0.514530	0.457393
0.593606	0.397266	0.412793	0.431204
0.534382	0.464741	0.458641	0.417299
0.521924	0.404541	0.392418	0.624609
0.571339	0.543937	0.343894	0.379259
0.628681	0.680485	0.396836	0.378522
0.587904	0.462116	0.326873	0.440864
0.600992	0.540494	0.417064	0.349167
0.480155	0.346121	0.602736	0.316015
0.503191	0.537891	0.593312	0.363699
0.572604	0.389360	0.404804	0.430824
0.534089	0.577297	0.599080	0.408154
0.554345	0.489568	0.514120	0.352823
0.560035	0.407987	0.252889	0.368411
0.604313	0.414195	0.566135	0.404395
0.574155	0.505573	0.424203	0.395749
0.570568	0.477283	0.219707	0.447135
0.493925	0.587282	0.593501	0.278440
0.607732	0.611498	0.540928	0.418678
0.569141	0.561094	0.553067	0.441914
0.560559	0.495731	0.386333	0.395447
0.624414	0.531289	0.301911	0.374005
0.632401	0.541135	0.448661	0.442877
0.585553	0.537106	0.513108	0.344947
0.556984	0.617248	0.667831	0.362820
0.520338	0.491704	0.210540	0.318166
0.522139	0.423068	0.545161	0.410346
0.556126	0.553643	0.660494	0.380295
0.524704	0.507274	0.650950	0.446071
0.505392	0.688899	0.546388	0.376950
0.488965	0.537929	0.572360	0.345153
0.541419	0.474365	0.634014	0.575410
0.495166	0.484491	0.498862	0.307387
0.579382	0.508451	0.460622	0.344674
0.542857	0.481824	0.385637	0.385117
0.609351	0.510396	0.440646	0.423635
0.525570	0.550105	0.418215	0.360521
0.554614	0.572657	0.401952	0.338906
0.551149	0.481490	0.392692	0.374623
0.557321	0.476740	0.406792	0.414472
0.593104	0.549101	0.430742	0.416586
0.511967	0.658690	0.386931	0.339964
0.558539	0.399696	0.568310	0.375470
0.519710	0.527100	0.469058	0.385331
0.563296	0.579664	0.422721	0.421097
0.549662	0.485171	0.494970	0.385258
0.527965	0.436297	0.241681	0.372544
0.565701	0.560034	0.733367	0.477279
0.563731	0.498434	0.209724	0.329020
0.575849	0.418204	0.520982	0.390257
0.578790	0.419531	0.386457	0.353079
0.570137	0.660870	0.731236	0.444461
0.544167	0.626064	0.295044	0.349507
0.525863	0.550049	0.644450	0.334648
0.600822	0.509487	0.654979	0.457482
0.555955	0.404606	0.466776	0.390157
0.565821	0.520103	0.549729	0.492489
0.534117	0.459643	0.545646	0.373238
0.698874	0.519265	0.544862	0.481119
0.506389	0.790262	0.457616	0.281971
0.586430	0.440464	0.524349	0.386866
0.564730	0.522523	0.387012	0.369622
0.451899	0.526390	0.592124	0.322081
0.556512	0.457018	0.253051	0.414886
0.608491	0.405867	0.405221	0.415781
0.558717	0.520725	0.432463	0.402661
0.507443	0.486107	0.710366	0.326942
0.590680	0.401430	0.353250	0.472570
0.569140	0.603802	0.542671	0.477538
0.560537	0.527750	0.481392	0.406185
0.647428	0.629767	0.365918	0.362047
0.550481	0.537540	0.479610	0.475301
0.502054	0.508076	0.331230	0.412566
0.572033	0.458005	0.158894	0.383438
0.474096	0.497083	0.449824	0.319237
0.458133	0.503370	0.386610	0.415273
0.540319	0.573741	0.478375	0.341585
0.566869	0.646777	0.646846	0.310636
0.457491	0.586812	0.582764	0.394147
0.555377	0.514684	0.380843	0.332182
0.490521	0.514998	0.473114	0.503080
0.563148	0.497894	0.427336	0.412938
0.525567	0.498645	0.500981	0.353692
0.579596	0.466666	0.335341	0.441261
0.599052	0.630852	0.482525	0.394749
0.532929	0.497762	0.431518	0.347832
0.555871	0.436469	0.579600	0.444695
0.544791	0.565292	0.561541	0.405939
0.522116	0.522881	0.459514	0.366005
0.592454	0.437790	0.432292	0.359087
0.605221	0.415054	0.350802	0.380092
0.607409	0.524001	0.387608	0.453868
0.535878	0.509733	0.326726	0.396450
0.575755	0.551890	0.341823	0.362073
0.608900	0.547716	0.569314	0.376473
0.527017	0.541159	0.578211	0.419317
0.535129	0.509911	0.409848	0.467585
0.542163	0.489338	0.304138	0.422431
0.561223	0.492660	0.467770	0.419296
0.572730	0.493334	0.561393	0.359086
0.595713	0.573896	0.537037	0.401083
0.491928	0.391156	0.771044	0.372092
0.498743	0.455395	0.655078	0.372951
0.559045	0.485956	0.592600	0.338588
0.502299	0.513169	0.372265	0.329785
0.609876	0.479793	0.552649	0.413503
0.466489	0.518687	0.357642	0.445671
0.519113	0.598488	0.555782	0.303972
0.511066	0.430728	0.404354	0.381744
0.665857	0.510662	0.408579	0.397807
0.551448	0.444160	0.563338	0.369755
0.519342	0.452295	0.600195	0.409428
0.498623	0.394853	0.296197	0.318769
0.554488	0.576374	0.289400	0.357675
0.533053	0.574060	0.371712	0.338418
0.508865	0.466735	0.380992	0.443725
0.564198	0.505363	0.377624	0.336451
0.578963	0.504184	0.381551	0.436794
0.562007	0.542190	0.389431	0.377868
0.552594	0.460700	0.706501	0.487112
0.530240	0.617003	0.271698	0.316912
0.499658	0.437666	0.665427	0.345625
0.600717	0.610829	0.447911	0.407148
0.552877	0.625569	0.634917	0.345773
0.556537	0.517300	0.595393	0.455266
0.493098	0.420205	0.394645	0.431901
0.558561	0.378381	0.487301	0.370257
0.622267	0.541232	0.426655	0.377820
0.599876	0.262775	0.578039	0.397777
0.517485	0.491923	0.596406	0.359808
0.604055	0.654860	0.487614	0.338530
0.562251	0.515955	0.309610	0.440540
0.607098	0.512912	0.555118	0.538029
0.519259	0.372946	0.396134	0.372035
0.601749	0.487082	0.555718	0.400614
0.551218	0.512837	0.172557	0.472196
0.527436	0.486252	0.386912	0.437837
0.558766	0.518881	0.422214	0.480533
0.601606	0.433845	0.461259	0.381237
0.540307	0.540905	0.312973	0.479234
0.553949	0.511514	0.317194	0.323664
0.634674	0.579763	0.519530	0.379287
0.519820	0.460692	0.574213	0.439772
0.590429	0.453514	0.562167	0.425192
0.519678	0.454654	0.282818	0.398959
0.564837	0.473498	0.547435	0.421466
0.526628	0.512980	0.373343	0.410556
0.586640	0.409118	0.292021	0.454170
0.526550	0.524337	0.153892	0.304987
0.486966	0.520179	0.333613	0.343127
0.507421	0.500725	0.355511	0.402650
0.545652	0.504126	0.297167	0.348568
0.543226	0.564712	0.501536	0.485995
0.551027	0.470558	0.531145	0.399702
0.594111	0.521423	0.235495	0.386367
0.547998	0.469505	0.582002	0.467376
0.516933	0.451108	0.458886	0.345640
0.559034	0.585327	0.350466	0.391828
0.546827	0.403454	0.120431	0.347510
0.510662	0.455614	0.283763	0.340890
0.533958	0.476182	0.495424	0.433341
0.592250	0.488106	0.495648	0.405867
0.498527	0.397774	0.333437	0.343550
0.613539	0.551436	0.527135	0.401972
0.578557	0.391697	0.283925	0.382609
0.578875	0.454054	0.625315	0.384648
0.495951	0.549760	0.430731	0.320174
0.593034	0.467054	0.444723	0.443847
0.589106	0.457468	0.653355	0.370528
0.549444	0.556465	0.335054	0.328695
0.653501	0.538941	0.367073	0.395655
0.519928	0.471081	0.451226	0.366144
0.579603	0.597510	0.310879	0.372933
0.583424	0.560315	0.324382	0.343674
0.615304	0.498153	0.427835	0.396297
0.523752	0.583648	0.350265	0.333511
0.561139	0.470825	0.313728	0.466759
0.571948	0.589479	0.552858	0.362329
0.593725	0.549007	0.710670	0.477972
0.599852	0.427411	0.208357	0.513524
0.596929	0.573113	0.339060	0.348981
0.541989	0.524170	0.347180	0.406176
0.503902	0.568606	0.488493	0.400357
0.493830	0.684566	0.212886	0.296145
0.515934	0.414772	0.683161	0.347297
0.526842	0.341139	0.409469	0.436358
0.616849	0.599087	0.382473	0.369336
0.584128	0.480570	0.545138	0.386592
0.506453	0.663786	0.390958	0.285638
0.579692	0.560492	0.412830	0.468508
0.600692	0.487557	0.405988	0.409838
0.567243	0.621747	0.339838	0.460033
0.535277	0.550207	0.270195	0.497832
0.546520	0.412877	0.302972	0.349165
0.515370	0.444779	0.453729	0.315441
0.525172	0.666619	0.408010	0.361076
0.613559	0.526346	0.508293	0.389052
0.542508	0.456497	0.649895	0.403877
0.507484	0.474491	0.550307	0.405414
0.525725	0.470735	0.690023	0.472363
0.537477	0.405022	0.361121	0.430057
0.503040	0.622484	0.455956	0.288501
0.570487	0.506297	0.420551	0.364190
0.551331	0.523401	0.453360	0.342355
0.602274	0.539345	0.481897	0.450790
0.546865	0.560651	0.424944	0.442425
0.506871	0.356330	0.418940	0.341785
0.547043	0.609686	0.350017	0.359996
0.567524	0.605264	0.878037	0.442318
0.548238	0.606691	0.664347	0.322823
0.573536	0.419435	0.562829	0.533707
0.584550	0.604159	0.496788	0.354634
0.553249	0.465668	0.509780	0.495683
0.584256	0.524961	0.449019	0.455105
0.518068	0.456456	0.661494	0.373794
0.494369	0.486111	0.348607	0.312925
0.585229	0.453025	0.422439	0.487236
0.523330	0.532865	0.232555	0.373021
0.656779	0.448454	0.273129	0.520304
0.581415	0.413986	0.470204	0.367750
0.612511	0.501299	0.495409	0.420933
0.553783	0.620189	0.197332	0.341818
0.607051	0.400681	0.337098	0.397122
0.538538	0.501618	0.451482	0.393357
0.563201	0.542549	0.589454	0.430702
0.550060	0.480739	0.571606	0.402192
0.616313	0.450918	0.481131	0.419234
0.598703	0.476473	0.415458	0.402408
0.562541	0.715025	0.386352	0.295900
0.585509	0.524265	0.318033	0.514455
0.501154	0.495151	0.820538	0.385017
0.531236	0.432147	0.411442	0.444340
0.537581	0.595852	0.438041	0.328825
0.544022	0.606069	0.493978	0.310676
0.476348	0.498642	0.265923	0.324888
0.620918	0.510241	0.285098	0.398399
0.506985	0.618078	0.353507	0.359348
0.566387	0.466629	0.382630	0.419516
0.536319	0.645059	0.464396	0.444638
0.594017	0.534912	0.493640	0.356450
0.548316	0.511476	0.522963	0.324385
0.551770	0.315911	0.248662	0.385643
0.650392	0.406223	0.545527	0.510584
0.615813	0.552908	0.460635	0.427799
0.533193	0.625247	0.617760	0.376075
0.596226	0.381791	0.442969	0.446457
0.527886	0.458456	0.486384	0.392417
0.564995	0.555009	0.454157	0.406982
0.610819	0.427016	0.516389	0.392146
0.547986	0.354244	0.236000	0.541880
0.541506	0.574945	0.583118	0.349565
0.567278	0.531096	0.222230	0.332308
0.547774	0.486658	0.269135	0.455912
0.534353	0.516555	0.679307	0.414927
0.573651	0.393822	0.233291	0.361795
0.562996	0.594452	0.543999	0.319319
0.655981	0.445460	0.380090	0.402748
0.526631	0.486840	0.422507	0.354357
0.712242	0.574013	0.354299	0.416451
0.556491	0.459885	0.432749	0.378562
0.597271	0.560328	0.169712	0.345290
0.638002	0.498625	0.279721	0.402039
0.528897	0.427470	0.392489	0.350737
0.561170	0.568102	0.340748	0.328872
0.593479	0.542730	0.274030	0.374671
0.506211	0.546492	0.844007	0.334013
0.496940	0.539534	0.891675	0.340120
0.619415	0.493277	0.440591	0.385759
0.562481	0.540763	0.606975	0.514270
0.556014	0.430403	0.583680	0.383588
0.436997	0.458623	0.381075	0.317383
0.591704	0.457188	0.362337	0.458980
0.552176	0.429246	0.455445	0.433922
0.572456	0.472663	0.453522	0.545982
0.558473	0.544769	0.354293	0.324299
0.498808	0.678103	0.465310	0.349009
0.551896	0.615571	0.344005	0.486124
0.593173	0.515327	0.383231	0.346595
0.509254	0.276932	0.257703	0.338049
0.599016	0.641399	0.113845	0.394987
0.601551	0.574752	0.413036	0.380883
0.493412	0.430212	0.527224	0.318737
0.557226	0.434694	0.330503	0.408940
0.567216	0.580506	0.250342	0.399066
0.464887	0.526467	0.518944	0.455392
0.560943	0.568591	0.519120	0.387924
0.567187	0.357417	0.469854	0.361383
0.514578	0.489254	0.282554	0.366111
0.569341	0.519953	0.537175	0.498171
0.460485	0.535181	0.634313	0.301980
0.569837	0.592772	0.393694	0.324219
0.572658	0.493067	0.213851	0.473512
0.597639	0.475841	0.450767	0.357619
0.611449	0.381747	0.436732	0.387283
0.610302	0.563369	0.306035	0.472068
0.556116	0.374755	0.541954	0.370916
0.659187	0.474392	0.375906	0.582200
0.568084	0.454688	0.427480	0.413428
0.579875	0.420442	0.493437	0.410837
0.570616	0.263359	0.277650	0.427328
0.647078	0.572520	0.256005	0.487565
0.551780	0.500516	0.592755	0.341882
0.521941	0.464970	0.395143	0.445730
0.611379	0.416102	0.519280	0.400993
0.490518	0.543934	0.377582	0.437865
0.531156	0.557353	0.389680	0.389848
0.635976	0.608853	0.717227	0.363179
0.555672	0.436873	0.671938	0.456640
0.512219	0.397040	0.517849	0.356749
0.668660	0.566676	0.496675	0.512365
0.526432	0.550483	0.598500	0.345565
0.502096	0.502672	0.488738	0.313546
0.571431	0.599392	0.340904	0.324958
0.567845	0.634993	0.527295	0.325716
0.571410	0.472287	0.358194	0.423235
0.501877	0.549534	0.446756	0.312750
0.587277	0.480949	0.531182	0.353450
0.590072	0.471590	0.690251	0.388942
0.600437	0.561355	0.454116	0.461041
0.497976	0.558120	0.658944	0.393667
0.563427	0.574705	0.139238	0.341957
0.509321	0.557906	0.520680	0.518149
0.518017	0.474520	0.382623	0.529847
0.506771	0.446559	0.195306	0.347570
0.468783	0.646114	0.367645	0.398168
0.571586	0.500971	0.399908	0.415789
0.540492	0.530895	0.618518	0.400932
0.592760	0.630432	0.493771	0.449302
0.535342	0.555672	0.442324	0.319614
0.499653	0.503266	0.394885	0.295803
0.487247	0.612018	0.537283	0.423025
0.529352	0.434576	0.585541	0.328028
0.466361	0.360996	0.411388	0.404892
0.478572	0.531720	0.479800	0.355950
0.515752	0.609146	0.479972	0.408180
0.559410	0.482515	0.397294	0.358220
0.500778	0.534849	0.412450	0.437236
0.668982	0.469428	0.513264	0.401407
0.513794	0.519284	0.380430	0.436589
0.568200	0.516660	0.528937	0.398834
0.574269	0.555999	0.496918	0.331194
0.559534	0.606470	0.670017	0.502838
0.536443	0.617050	0.650547	0.334880
0.561679	0.584720	0.490014	0.516741
0.533596	0.550979	0.468252	0.309758
0.509577	0.411332	0.499895	0.363961
0.515907	0.558504	0.252443	0.324997
0.535221	0.460841	0.495005	0.375373
0.581182	0.471462	0.268868	0.346649
0.513661	0.588769	0.250653	0.296462
0.616486	0.522285	0.398759	0.397511
0.570534	0.537387	0.285832	0.375446
0.544530	0.433024	0.572800	0.458320
0.637468	0.468618	0.574325	0.418328
0.572098	0.464509	0.394971	0.342937
0.540634	0.497762	0.386587	0.377673
0.554760	0.468369	0.294149	0.402079
0.613235	0.450352	0.443059	0.388873
0.608413	0.405165	0.597674	0.442832
0.605104	0.545142	0.319910	0.366047
0.554737	0.577566	0.488707	0.495907
0.560422	0.484235	0.394141	0.381281
0.555762	0.576417	0.481134	0.489243
0.644932	0.590964	0.521177	0.405402
0.542781	0.460571	0.620418	0.341685
0.506002	0.441837	0.677663	0.555314
0.457100	0.620834	0.466961	0.380070
0.528922	0.596777	0.369027	0.356204
0.604477	0.493598	0.562021	0.423983
0.501355	0.555882	0.309918	0.317808
0.556531	0.328648	0.388158	0.416079
0.502662	0.511727	0.285122	0.301875
0.603558	0.581172	0.337643	0.348609
0.523377	0.442118	0.526279	0.377481
0.638043	0.356569	0.298124	0.441186
0.544283	0.484106	0.273950	0.422249
0.521717	0.459253	0.413171	0.403057
0.550092	0.534231	0.538954	0.442789
0.463300	0.507132	0.358330	0.381279
0.720558	0.514411	0.672566	0.441643
0.522123	0.523294	0.373500	0.342664
0.625070	0.512156	0.415089	0.439219
0.535383	0.420052	0.287254	0.355064
0.667264	0.477599	0.791932	0.436731
0.575591	0.513315	0.682290	0.375426
0.604873	0.382473	0.426923	0.442575
0.528119	0.534362	0.651109	0.416767
0.571807	0.543926	0.333936	0.509524
0.561891	0.509562	0.559624	0.367535
0.658144	0.614150	0.458833	0.377935
0.536837	0.589696	0.594899	0.313203
0.616485	0.556291	0.276753	0.380049
0.530913	0.656602	0.540997	0.324719
0.551677	0.590979	0.558063	0.317064
0.577934	0.647688	0.435853	0.319634
0.526620	0.473809	0.358400	0.398756
0.519624	0.427230	0.444335	0.333868
0.546372	0.699090	0.322622	0.295601
0.616289	0.595390	0.285483	0.463357
0.651494	0.493147	0.564802	0.532641
0.589997	0.466214	0.455138	0.363985
0.571536	0.554964	0.714881	0.334044
0.564737	0.524849	0.316914	0.368375
0.566852	0.715861	0.498183	0.394287
0.611709	0.588074	0.703426	0.463508
0.485966	0.497086	0.360169	0.326149
0.544752	0.426680	0.448118	0.352021
0.607515	0.571132	0.140809	0.355352
0.605663	0.626367	0.478063	0.366651
0.595724	0.656876	0.447409	0.335471
0.579437	0.444904	0.432143	0.384377
0.579268	0.467248	0.455430	0.423220
0.488249	0.481118	0.426981	0.410845
0.536309	0.485097	0.306818	0.354989
0.552244	0.608412	0.391462	0.380234
0.504196	0.448786	0.527501	0.364996
0.497925	0.460381	0.410128	0.340096
0.594451	0.679140	0.265238	0.403557
0.582125	0.510376	0.221093	0.358915
0.595798	0.542806	0.626359	0.426328
0.518147	0.489984	0.440576	0.361179
0.542001	0.392002	0.501830	0.499650
0.508872	0.493658	0.575345	0.385642
0.613572	0.578354	0.373684	0.366599
0.543927	0.461211	0.549179	0.367663
0.545942	0.518357	0.472515	0.386814
0.613795	0.462082	0.471319	0.420871
0.504948	0.473506	0.536802	0.413285
0.608479	0.493651	0.356835	0.407604
0.622548	0.624712	0.455572	0.363164
0.538874	0.522682	0.440427	0.362160
0.628234	0.533077	0.203510	0.499779
0.507642	0.576874	0.494454	0.300536
0.521873	0.569372	0.462046	0.464275
0.578537	0.423170	0.499650	0.383861
0.596114	0.493111	0.619446	0.389219
0.600105	0.552455	0.491538	0.349607
0.573636	0.625500	0.358050	0.393216
0.622954	0.534677	0.334167	0.380698
0.559522	0.615748	0.445424	0.312379
0.595749	0.409837	0.441755	0.400226
0.597014	0.516121	0.551591	0.378575
0.599419	0.455797	0.241403	0.359211
0.505821	0.521898	0.585286	0.433608
0.548502	0.451550	0.697827	0.354435
0.558941	0.514544	0.538271	0.357040
0.600153	0.463195	0.559465	0.389559
0.602160	0.441721	0.460282	0.380235
0.588407	0.554166	0.392059	0.398804
0.685967	0.493188	0.291478	0.422105
0.547422	0.564667	0.606208	0.429537
0.534757	0.496059	0.436199	0.422972
0.573136	0.403564	0.558713	0.363891
0.540664	0.445479	0.370696	0.417058
0.637725	0.570199	0.293455	0.365669
0.636858	0.439346	0.696109	0.412222
0.564400	0.493544	0.343201	0.377591
0.589029	0.486423	0.649761	0.352967
0.545958	0.489647	0.561710	0.350252
0.582283	0.415417	0.190338	0.365013
0.610324	0.607383	0.500090	0.344704
0.467264	0.516290	0.697306	0.380482
0.537837	0.439729	0.390169	0.338225
0.523821	0.621663	0.711917	0.342733
0.579460	0.473778	0.238632	0.458328
0.574512	0.575903	0.528945	0.339208
0.568532	0.497083	0.454118	0.375183
0.638665	0.412987	0.364961	0.469997
0.532758	0.613881	0.585711	0.416740
0.527773	0.565938	0.339992	0.445880
0.489835	0.420901	0.365151	0.447420
0.555009	0.668001	0.511947	0.521176
0.579767	0.643315	0.319217	0.374822
0.531831	0.585358	0.324917	0.384869
0.617926	0.601930	0.422244	0.363206
0.549662	0.497579	0.547789	0.411062
0.505140	0.470769	0.290876	0.395552
0.553774	0.504718	0.416659	0.349245
0.513880	0.532345	0.403144	0.308221
0.613894	0.461778	0.266708	0.393509
0.523794	0.652429	0.370624	0.333202
0.482332	0.536217	0.735084	0.400180
0.581698	0.503430	0.318035	0.398433
0.536664	0.580034	0.491424	0.315071
0.668125	0.544769	0.550114	0.404284
0.544890	0.601358	0.313503	0.326331
0.607124	0.494455	0.639317	0.450639
0.504360	0.533563	0.415901	0.448010
0.526992	0.437302	0.500373	0.420919
0.709098	0.599454	0.314012	0.473356
0.590015	0.649886	0.399563	0.334123
0.571315	0.570436	0.553736	0.347625
0.526876	0.413789	0.461786	0.327074
0.602506	0.489667	0.499255	0.368890
0.547479	0.614407	0.428643	0.363891
0.495730	0.460399	0.485989	0.300308
0.551698	0.463098	0.489860	0.339257
0.598248	0.567098	0.390078	0.441042
0.484114	0.557749	0.436745	0.323071
0.561634	0.459350	0.483255	0.472799
0.602630	0.559117	0.587800	0.374852
0.550355	0.521222	0.540755	0.359543
0.561188	0.545702	0.578146	0.387527
0.537144	0.550893	0.597186	0.363431
0.562892	0.594080	0.311438	0.378332
0.626603	0.566723	0.581790	0.416999
0.590593	0.408425	0.231156	0.364815
0.607304	0.512327	0.393799	0.410787
0.570660	0.526095	0.378603	0.383747
0.562056	0.527775	0.246466	0.505616
0.538254	0.647215	0.365642	0.331230
0.630508	0.551368	0.526418	0.410573
0.540186	0.525589	0.395751	0.329402
0.595707	0.462233	0.493455	0.494108
0.530440	0.587593	0.592850	0.365471
0.549144	0.530043	0.525251	0.382383
0.556887	0.395531	0.552591	0.370120
0.552220	0.497432	0.427762	0.384391
0.568298	0.539641	0.625313	0.376692
0.562278	0.482913	0.686851	0.431439
0.628051	0.544696	0.526708	0.387904
0.506874	0.410547	0.704865	0.380485
0.558780	0.451308	0.367788	0.351098
0.516506	0.501093	0.443571	0.305438
0.608587	0.572591	0.220294	0.369439
0.480773	0.516414	0.319709	0.288865
0.517538	0.491699	0.484135	0.381268
0.542398	0.494306	0.441430	0.407357
0.599983	0.541093	0.556583	0.375409
0.583761	0.618748	0.344401	0.358812
0.564711	0.565955	0.458773	0.337810
0.566583	0.453080	0.633927	0.345444
0.588693	0.660374	0.360757	0.328310
0.531667	0.453510	0.316822	0.404862
0.553113	0.547151	0.312980	0.332667
0.563279	0.600908	0.637300	0.440819
0.603900	0.562624	0.352484	0.433553
0.577319	0.528689	0.275297	0.334552
0.557920	0.545519	0.418920	0.510410
0.579760	0.524760	0.145740	0.356868
0.510629	0.574135	0.515577	0.361351
0.618650	0.633972	0.743059	0.375058
0.504693	0.485914	0.572756	0.379960
0.522679	0.576500	0.649573	0.524253
0.495706	0.399961	0.413790	0.350239
0.538674	0.289546	0.565195	0.395651
0.547882	0.489153	0.529997	0.471265
0.539856	0.346845	0.251996	0.369252
0.526123	0.653228	0.581194	0.297020
0.498762	0.637158	0.549342	0.370831
0.635977	0.644682	0.498392	0.358030
0.537804	0.442130	0.310111	0.405980
0.543390	0.547053	0.209247	0.325203
0.634707	0.510789	0.607098	0.496167
0.596035	0.496110	0.271148	0.429341
0.533808	0.660245	0.612753	0.288120
0.609348	0.543883	0.310481	0.387947
0.499994	0.549053	0.403328	0.383321
0.583588	0.554844	0.458912	0.458504
0.589261	0.542571	0.181581	0.432396
0.511014	0.392841	0.574926	0.531871
0.603668	0.483257	0.479498	0.439997
0.555189	0.623166	0.228431	0.419666
0.578284	0.531147	0.508960	0.399578
0.574320	0.496998	0.549761	0.400661
0.526543	0.488314	0.113716	0.317608
0.577389	0.545754	0.401751	0.473438
0.523380	0.361451	0.567260	0.351725
0.452977	0.423240	0.410778	0.383021
0.525778	0.464783	0.470554	0.337960
0.557990	0.521410	0.720940	0.358491
0.588959	0.325779	0.719199	0.397997
0.601980	0.409755	0.533049	0.427546
0.517393	0.526127	0.901582	0.336096
0.679988	0.474158	0.608251	0.453782
0.570336	0.497526	0.511533	0.498610
0.605474	0.593330	0.406031	0.434413
0.576721	0.439770	0.301165	0.564156
0.451013	0.605180	0.348301	0.303458
0.582963	0.513973	0.465142	0.490032
0.560296	0.460303	0.376300	0.415974
0.584681	0.585281	0.419287	0.365484
0.619026	0.578717	0.168214	0.405805
0.535462	0.443841	0.295532	0.333397
0.549762	0.449372	0.498747	0.382809
0.524998	0.448122	0.438523	0.357247
0.569778	0.514075	0.386490	0.423882
0.505898	0.499612	0.401854	0.381081
0.537926	0.453724	0.568150	0.429221
0.581609	0.508132	0.438647	0.465706
0.589613	0.616539	0.427992	0.398774
0.550010	0.573273	0.526729	0.490991
0.555861	0.516737	0.522883	0.433081
0.569227	0.610991	0.402995	0.387157
0.549575	0.460227	0.565039	0.344190
0.557302	0.541463	0.402042	0.444521
0.596917	0.622670	0.566475	0.452947
0.557301	0.557964	0.679824	0.342030
0.526618	0.562565	0.333848	0.516933
0.544483	0.547087	0.544532	0.385360
0.556529	0.538713	0.332185	0.336885
0.587934	0.512601	0.247082	0.342851
0.614406	0.470764	0.421998	0.435106
0.520243	0.410021	0.236937	0.338670
0.510833	0.487160	0.625021	0.425171
0.575544	0.471239	0.543277	0.448815
0.528747	0.564258	0.393497	0.384898
0.465102	0.503382	0.373907	0.458807
0.482518	0.481168	0.365152	0.293504
0.549829	0.586355	0.520186	0.311335
0.534946	0.478878	0.260435	0.385723
0.582006	0.517195	0.227631	0.475911
0.612689	0.612426	0.421693	0.447728
0.595400	0.445404	0.324992	0.375469
0.529887	0.456149	0.743836	0.363350
0.557415	0.586390	0.085244	0.370728
0.598259	0.518757	0.292342	0.389126
0.608961	0.451347	0.300502	0.367136
0.544761	0.509686	0.194291	0.477535
0.599223	0.522985	0.500323	0.360466
0.527731	0.371756	0.378154	0.372484
0.614050	0.512251	0.612182	0.401436
0.504868	0.455546	0.712360	0.365049
0.534205	0.568000	0.439467	0.321143
0.552257	0.616739	0.427604	0.446101
0.523842	0.525306	0.325357	0.334882
0.545550	0.542188	0.343511	0.382708
0.567745	0.570743	0.528578	0.409962
0.547616	0.574053	0.598733	0.418429
0.603411	0.538050	0.422872	0.386018
0.527667	0.538643	0.308118	0.442713
0.525193	0.560536	0.751097	0.345663
0.544623	0.546738	0.182116	0.314328
0.514925	0.422391	0.558247	0.415350
0.474063	0.556409	0.431644	0.307819
0.608960	0.541475	0.378634	0.435860
0.479420	0.394906	0.498620	0.348829
0.548571	0.476673	0.438066	0.348494
0.577290	0.345775	0.250579	0.478324
0.571478	0.497102	0.539419	0.340237
0.488606	0.537393	0.491211	0.335662
0.586497	0.562800	0.089603	0.334584
0.623709	0.572612	0.392174	0.438008
0.548830	0.448119	0.573213	0.364719
0.558418	0.224979	0.540130	0.418875
0.558858	0.401500	0.344714	0.478550
0.545805	0.509054	0.528611	0.337756
0.577995	0.419674	0.471973	0.361490
0.633109	0.412281	0.548126	0.422102
0.591083	0.523401	0.466888	0.417757
0.642204	0.624435	0.470112	0.424181
0.599561	0.607187	0.543184	0.406162
0.507978	0.550997	0.274833	0.347474
0.554952	0.699252	0.717971	0.438622
0.510262	0.485616	0.281045	0.393330
0.558914	0.401767	0.789134	0.357807
0.551842	0.615352	0.462958	0.319386
0.487530	0.572895	0.289187	0.378698
0.645346	0.591930	0.443909	0.424942
0.555091	0.421550	0.585652	0.378659
0.520006	0.436826	0.619866	0.373567
0.570014	0.261657	0.750203	0.485032
0.543999	0.507730	0.609827	0.388291
0.591339	0.467234	0.559011	0.398832
0.576617	0.576431	0.316184	0.343066
0.555859	0.551629	0.391218	0.488837
0.607972	0.581175	0.524243	0.413257
0.541909	0.497722	0.430583	0.327107
0.541195	0.471989	0.387465	0.333808
0.525137	0.528986	0.285560	0.466408
0.571394	0.557719	0.375979	0.389078
0.566848	0.475532	0.455593	0.364456
0.579806	0.427970	0.492749	0.357521
0.623113	0.595269	0.565994	0.420947
0.572613	0.545658	0.585529	0.402574
0.530056	0.462050	0.538616	0.341755
0.540066	0.488229	0.261497	0.352788
0.566419	0.587286	0.503171	0.349963
0.567293	0.318970	0.404966	0.457147
0.545598	0.506746	0.378415	0.340269
0.507258	0.372395	0.355451	0.403878
0.536918	0.451063	0.560445	0.391109
0.496696	0.507490	0.507421	0.361528
0.502249	0.564189	0.395267	0.364863
0.594516	0.501368	0.431700	0.403145
0.626018	0.494941	0.542523	0.385701
0.665823	0.545923	0.255780	0.455623
0.602237	0.447460	0.380804	0.506921
0.539634	0.494937	0.462871	0.386784
0.536785	0.582355	0.647590	0.324038
0.500125	0.557718	0.354596	0.441148
0.514936	0.493669	0.449457	0.515678
0.609185	0.331311	0.479201	0.422175
0.562362	0.474189	0.314854	0.436617
0.477309	0.394342	0.437257	0.443226
0.494864	0.350868	0.306988	0.328268
0.520654	0.386742	0.480708	0.384574
0.630484	0.393999	0.591777	0.469142
0.515746	0.516495	0.269845	0.324214
0.562782	0.436664	0.570439	0.392278
0.501888	0.591484	0.566855	0.308877
0.492934	0.480843	0.505779	0.339282
0.557738	0.500479	0.514759	0.348216
0.547353	0.556326	0.404074	0.361294
0.522398	0.654969	0.617748	0.331955
0.526757	0.609282	0.367263	0.367035
0.568842	0.545857	0.327412	0.516415
0.471683	0.568520	0.430841	0.369433
0.499516	0.500465	0.529172	0.342876
0.593386	0.408704	0.472906	0.462256
0.543292	0.671256	0.601452	0.323378
0.536396	0.532850	0.321355	0.343528
0.500089	0.420533	0.500959	0.450958
0.585511	0.490243	0.658906	0.384617
0.577724	0.436958	0.331635	0.412046
0.568696	0.481197	0.652034	0.497882
0.617577	0.666063	0.422969	0.400803
0.558980	0.493603	0.587368	0.345512
0.595779	0.521631	0.288550	0.489401
0.541747	0.565448	0.453465	0.360752
0.548289	0.648126	0.566266	0.368585
0.619716	0.419034	0.382060	0.408400
0.626721	0.584055	0.378586	0.365672
0.530669	0.580911	0.296122	0.366296
0.568499	0.498772	0.411238	0.535374
0.582112	0.560779	0.327761	0.343665
0.554497	0.402641	0.242513	0.369861
0.558974	0.500647	0.532288	0.516137
0.645805	0.546527	0.519559	0.416591
0.536877	0.502380	0.349389	0.408806
0.528462	0.585527	0.308591	0.299502
0.626118	0.525999	0.500584	0.382054
0.491967	0.497873	0.273145	0.364506
0.507142	0.402732	0.108732	0.326976
0.616132	0.456315	0.317031	0.425104
0.616607	0.540226	0.819304	0.373222
0.497971	0.469809	0.326015	0.346130
0.567487	0.465457	0.369453	0.443230
0.553563	0.601943	0.480487	0.327233
0.531424	0.393272	0.443772	0.374713
0.497339	0.414615	0.651640	0.323804
0.500217	0.523949	0.685314	0.312135
0.544988	0.482581	0.330183	0.331949
0.595841	0.469237	0.506576	0.376765
0.530533	0.490347	0.498676	0.408981
0.498143	0.583167	0.703152	0.455251
0.602269	0.518017	0.490538	0.388677
0.540659	0.608785	0.365881	0.337748
0.592911	0.459924	0.536302	0.394337
0.562169	0.591733	0.342408	0.342653
0.579110	0.598818	0.545427	0.433288
0.640221	0.522340	0.423179	0.440137
0.523734	0.510342	0.807395	0.369459
0.629062	0.467410	0.414042	0.384502
0.533226	0.502444	0.504456	0.324896
0.612198	0.518541	0.543750	0.363741
0.566165	0.537423	0.192457	0.339475
0.579569	0.556033	0.570402	0.384166
0.537624	0.623899	0.524423	0.361025
0.611363	0.477335	0.365006	0.390334
0.635646	0.598473	0.411836	0.423507
0.614532	0.430388	0.653388	0.431368
0.645776	0.514379	0.418977	0.391820
0.596943	0.347425	0.416815	0.381678
0.479787	0.481943	0.387058	0.326795
0.545786	0.678580	0.399871	0.342692
0.520521	0.582825	0.133080	0.426551
0.551098	0.514721	0.244793	0.438212
0.598200	0.466182	0.706141	0.450620
0.558620	0.483256	0.630576	0.348297
0.519487	0.492258	0.501861	0.371763
0.474920	0.614621	0.413845	0.356248
0.499217	0.396901	0.512141	0.330444
0.601641	0.486868	0.533575	0.364618
0.515855	0.405843	0.394081	0.332478
0.584265	0.540079	0.565789	0.369576
0.544643	0.448385	0.264394	0.332228
0.552935	0.577466	0.476487	0.501735
0.483130	0.408120	0.508590	0.371558
0.613968	0.508495	0.333704	0.378716
0.554232	0.469747	0.263193	0.382494
0.558164	0.516321	0.574342	0.331058
0.577694	0.484114	0.374218	0.369538
0.552949	0.545869	0.315300	0.390515
0.561405	0.472829	0.432777	0.646400
0.570946	0.444524	0.411960	0.369873
0.578235	0.634657	0.515313	0.340832
0.506714	0.548681	0.464591	0.290928
0.493726	0.448402	0.516735	0.348837
0.545287	0.430371	0.427415	0.341953
0.592433	0.625632	0.477389	0.340545
0.662145	0.468393	0.434037	0.413232
0.530338	0.555654	0.632638	0.366028
0.526523	0.663001	0.400481	0.431014
0.537078	0.569508	0.301500	0.384521
0.552434	0.573166	0.593580	0.354843
0.559553	0.495938	0.530861	0.343533
0.537277	0.566891	0.636439	0.372194
0.435299	0.460671	0.167223	0.293266
0.548739	0.495291	0.463249	0.352885
0.622500	0.444714	0.570449	0.437425
0.562754	0.663375	0.489834	0.333753
0.571023	0.458770	0.263695	0.445700
0.490660	0.451473	0.508514	0.382659
0.506688	0.436275	0.388717	0.380867
0.440161	0.523675	0.536931	0.418206
0.645507	0.636615	0.584660	0.415057
0.583996	0.507760	0.363026	0.488910
0.556247	0.570006	0.662876	0.575886
0.552810	0.414800	0.377129	0.438653
0.635940	0.534972	0.384573	0.442317
0.580979	0.462679	0.167318	0.350585
0.564258	0.493532	0.381542	0.338275
0.568262	0.478309	0.469454	0.423101
0.578874	0.454218	0.392296	0.409738
0.571315	0.411594	0.276228	0.357549
0.534894	0.435192	0.293208	0.371471
0.622873	0.453670	0.517582	0.387148
0.583019	0.559477	0.432369	0.424748
0.520663	0.612186	0.569227	0.319125
0.581965	0.491298	0.365830	0.384945
0.610589	0.534628	0.569749	0.356646
0.602880	0.529139	0.592055	0.370509
0.512256	0.358267	0.606892	0.327557
0.567435	0.541396	0.347941	0.387030
0.566431	0.425058	0.570964	0.438399
0.580326	0.469796	0.482930	0.398067
0.628625	0.491888	0.431006	0.394518
0.553352	0.557432	0.413111	0.579660
0.568374	0.478115	0.464993	0.365719
0.563172	0.505067	0.207478	0.452913
0.491907	0.506464	0.548019	0.322507
0.518788	0.525829	0.486501	0.384542
0.520918	0.517133	0.364046	0.320529
0.569846	0.520347	0.382683	0.530776
0.540970	0.496826	0.387556	0.393364
0.548817	0.581733	0.776403	0.338908
0.576782	0.452452	0.355914	0.459423
0.621810	0.613264	0.499050	0.359501
0.517290	0.520134	0.407963	0.415740
0.545219	0.420340	0.462799	0.416726
0.547910	0.544176	0.511952	0.335188
0.588062	0.473187	0.472276	0.393288
0.593725	0.538685	0.449028	0.376702
0.550107	0.474327	0.357606	0.472582
0.553384	0.399654	0.706867	0.469942
0.581663	0.573040	0.000000	0.387797
0.540237	0.506617	0.228569	0.441743
0.551596	0.466452	0.442780	0.345488
0.543725	0.554883	0.491970	0.325390
0.669615	0.492307	0.611962	0.455553
0.542599	0.397477	0.588720	0.386455
0.490938	0.464996	0.613768	0.315741
0.493235	0.547359	0.672243	0.315829
0.518505	0.520624	0.514572	0.390951
0.547833	0.572578	0.115279	0.325854
0.546385	0.445259	0.642890	0.501006
0.592118	0.567718	0.492419	0.342033
0.530657	0.475831	0.233004	0.352467
0.542589	0.529060	0.239963	0.386510
0.556211	0.671651	0.372102	0.395358
0.534411	0.600770	0.508188	0.331601
0.525820	0.465882	0.440106	0.349253
0.588151	0.454506	0.324926	0.447773
0.488036	0.531236	0.582968	0.297175
0.531361	0.611300	0.450255	0.368789
0.553794	0.590550	0.476745	0.359929
0.705943	0.484780	0.603585	0.508402
0.534877	0.430946	0.294662	0.463437
0.565132	0.460822	0.685549	0.409212
0.581981	0.619706	0.419190	0.387208
0.537819	0.489645	0.562246	0.446721
0.572187	0.651772	0.460751	0.526361
0.522083	0.500714	0.362879	0.325779
0.567380	0.496270	0.527309	0.374881
0.592992	0.619960	0.457431	0.338148
0.579725	0.609299	0.097657	0.370650
0.569398	0.479448	0.304801	0.346547
0.614072	0.468520	0.386773	0.440638
0.581360	0.402711	0.389148	0.357845
0.516115	0.487830	0.320682	0.379239
0.606275	0.590726	0.426499	0.362860
0.551420	0.518997	0.356957	0.347934
0.548163	0.489498	0.292847	0.466807
0.502704	0.384935	0.378509	0.370035
0.491512	0.591585	0.766168	0.328899
0.581972	0.464327	0.514253	0.422554
0.597853	0.459671	0.533820	0.467471
0.588850	0.454805	0.533979	0.385099
0.518962	0.495202	0.455532	0.417209
0.545507	0.435211	0.463145	0.520049
0.570186	0.585608	0.611133	0.364974
0.574145	0.613891	0.728385	0.393555
0.587068	0.529469	0.362936	0.347089
0.474691	0.606624	0.323647	0.295885
0.586710	0.466940	0.377995	0.371532
0.612502	0.644115	0.284081	0.362758
0.511219	0.492032	0.288460	0.325693
0.548906	0.381194	0.605028	0.391077
0.572702	0.581250	0.244833	0.414442
0.525082	0.465652	0.343921	0.382707
0.562433	0.456409	0.303786	0.397218
0.556218	0.494847	0.540628	0.338445
0.594531	0.466260	0.134920	0.372604
0.526716	0.452385	0.410642	0.396880
0.635312	0.523518	0.441997	0.394620
0.524716	0.515981	0.643928	0.372907
0.547585	0.415333	0.220055	0.353525
0.546803	0.460382	0.556755	0.426442
0.641137	0.392268	0.672576	0.434398
0.566249	0.505956	0.127466	0.335245
0.540615	0.318128	0.395509	0.369640
0.535385	0.512702	0.386591	0.396692
0.605661	0.495667	0.266768	0.363081
0.628375	0.399742	0.567742	0.498735
0.599196	0.445248	0.385683	0.407540
0.609898	0.588863	0.417406	0.398368
0.586494	0.419998	0.633876	0.384628
0.535055	0.550545	0.512448	0.308421
0.519481	0.491186	0.256911	0.313678
0.514127	0.549969	0.503371	0.295513
0.597546	0.501419	0.404223	0.362690
0.613689	0.521894	0.542484	0.362442
0.475667	0.524185	0.270028	0.414145
0.534722	0.505664	0.320690	0.391860
0.622571	0.595483	0.315457	0.398427
0.514396	0.530044	0.612955	0.485703
0.555676	0.499484	0.517306	0.404419
0.608141	0.485997	0.376033	0.401117
0.524246	0.414304	0.688691	0.422354
0.575567	0.563134	0.406311	0.405232
0.536987	0.535925	0.618209	0.478661
0.537672	0.584259	0.358879	0.372113
0.526528	0.514565	0.437551	0.334067
0.535518	0.477354	0.347030	0.371629
0.567743	0.491010	0.515352	0.404476
0.553298	0.487633	0.528840	0.401027
0.572789	0.473702	0.530575	0.511389
0.554349	0.578058	0.544502	0.324378
0.529547	0.521040	0.435735	0.437088
0.557329	0.492795	0.316992	0.480157
0.538163	0.575052	0.383363	0.347236
0.561358	0.414477	0.293252	0.371496
0.530353	0.580305	0.232045	0.295164
0.634567	0.471168	0.546147	0.425253
0.464867	0.509819	0.417807	0.317302
0.504349	0.571680	0.465390	0.343269
0.553322	0.549664	0.514460	0.371336
0.490493	0.458096	0.270863	0.347010
0.513002	0.430962	0.157263	0.329775
0.577077	0.401112	0.496779	0.365074
0.487594	0.428266	0.236435	0.332246
0.561401	0.545121	0.229989	0.345189
0.548853	0.593270	0.255376	0.358100
0.537397	0.436212	0.723029	0.416414
0.496285	0.539387	0.395730	0.363585
0.576522	0.543691	0.416762	0.395702
0.502270	0.465323	0.569158	0.335207
0.600066	0.520896	0.433114	0.402341
0.609351	0.629915	0.265482	0.397384
0.559690	0.638173	0.676053	0.364945
0.488307	0.496447	0.334458	0.343371
0.614452	0.567630	0.692517	0.430234
0.531107	0.456090	0.525322	0.330589
0.587259	0.587761	0.163888	0.502959
0.536440	0.570717	0.412942	0.371484
0.582857	0.460287	0.261334	0.388003
0.563623	0.508226	0.621509	0.405095
0.474166	0.500184	0.388241	0.367807
0.532244	0.539514	0.545095	0.306968
0.509431	0.385686	0.518227	0.353515
0.650380	0.607464	0.575001	0.449410
0.613013	0.498731	0.509265	0.410441
0.547372	0.516781	0.278860	0.325825
0.571626	0.543842	0.493595	0.424092
0.469218	0.692412	0.610132	0.408920
0.677366	0.672484	0.665004	0.386486
0.625532	0.538740	0.437589	0.412466
0.620290	0.514665	0.380711	0.368484
0.501173	0.541083	0.409036	0.548684
0.650474	0.649966	0.295565	0.358222
0.547928	0.503718	0.409253	0.444781
0.563118	0.535052	0.544775	0.415067
0.608382	0.437598	0.407238	0.530333
0.507873	0.391493	0.452963	0.343024
0.500581	0.489498	0.604202	0.321674
0.512192	0.552232	0.316312	0.334213
0.542488	0.537781	0.704813	0.398027
0.455124	0.458680	0.372436	0.311980
0.464817	0.418461	0.502441	0.367127
0.562244	0.534418	0.783254	0.490701
0.492971	0.608594	0.403416	0.383445
0.553597	0.533511	0.538183	0.379799
0.528957	0.450705	0.708699	0.371693
0.575185	0.567656	0.403345	0.399706
0.474031	0.582398	0.528707	0.310237
0.590203	0.382538	0.449138	0.489278
0.489859	0.486766	0.376365	0.387258
0.501032	0.453841	0.395883	0.443075
0.509428	0.700576	0.449994	0.413959
0.508223	0.450631	0.411209	0.317271
0.548461	0.647351	0.506781	0.360819
0.518878	0.556122	0.338868	0.311074
0.495942	0.441003	0.361379	0.450359
0.590302	0.522807	0.377359	0.419174
0.538285	0.637662	0.360641	0.300605
0.541709	0.551402	0.452005	0.359510
0.462578	0.419325	0.227795	0.361755
0.620869	0.393481	0.312085	0.454098
0.517873	0.545252	0.414926	0.396576
0.522525	0.563913	0.610227	0.429491
0.585847	0.507775	0.601943	0.386829
0.549556	0.486169	0.384284	0.422513
0.534300	0.547504	0.341322	0.317077
0.504539	0.439655	0.617659	0.466266
0.486226	0.596877	0.705743	0.412439
0.590371	0.591181	0.359010	0.391002
0.569758	0.527154	0.374143	0.337032
0.500892	0.562398	0.304957	0.394332
0.517380	0.538559	0.577696	0.432831
0.562188	0.431069	0.244146	0.456636
0.531248	0.420656	0.732081	0.384750
0.575796	0.639300	0.503976	0.363424
0.542352	0.426129	0.323168	0.359777
0.557692	0.348178	0.349464	0.438595
0.618223	0.689177	0.364616	0.363464
0.581164	0.516053	0.652492	0.391295
0.538651	0.634182	0.459472	0.327829
0.575302	0.604707	0.207682	0.348399
0.572554	0.658286	0.554601	0.318982
0.536887	0.370299	0.361298	0.431159
0.567794	0.507504	0.311260	0.387650
0.496479	0.560569	0.406201	0.362775
0.599404	0.648755	0.541215	0.373170
0.606907	0.556120	0.565542	0.388322
0.545361	0.542235	0.400639	0.336806
0.616105	0.533769	0.440027	0.438051
0.710891	0.617796	0.554717	0.485828
0.568574	0.618584	0.531328	0.342209
0.566044	0.432534	0.556269	0.398606
0.522104	0.478236	0.517400	0.355579
0.636386	0.530233	0.372791	0.493957
0.650841	0.516988	0.339402	0.449409
0.641451	0.600043	0.418809	0.403084
0.618540	0.375514	0.382016	0.394060
0.550490	0.467609	0.526078	0.331292
0.520535	0.542894	0.515690	0.333269
0.605094	0.440149	0.654215	0.429800
0.612581	0.396056	0.705831	0.457208
0.570022	0.425024	0.275482	0.418944
0.554783	0.586649	0.512144	0.323972
0.527148	0.400089	0.370184	0.354208
0.600246	0.469291	0.634495	0.403584
0.550613	0.495100	0.508525	0.392478
0.532085	0.273866	0.391426	0.441705
0.634576	0.581266	0.211173	0.388911
0.584394	0.448831	0.467590	0.358990
0.610760	0.532698	0.475970	0.576293
0.590350	0.412345	0.251228	0.383537
0.561549	0.490793	0.376419	0.348161
0.547979	0.568849	0.595090	0.410722
0.516938	0.579613	0.357823	0.347975
0.597496	0.537017	0.346936	0.415748
0.563038	0.407169	0.342470	0.402110
0.520769	0.523834	1.000000	0.437191
0.537862	0.376932	0.496874	0.420731
0.526744	0.500394	0.376839	0.375607
0.522535	0.366561	0.416559	0.410478
0.584439	0.582697	0.576403	0.418480
0.633594	0.533232	0.582911	0.456606
0.579511	0.522833	0.280150	0.350938
0.484814	0.418599	0.525359	0.429860
0.574415	0.484933	0.507720	0.393094
0.514049	0.547261	0.416439	0.362413
0.553062	0.675011	0.559584	0.412677
0.574041	0.463831	0.604307	0.402826
0.607240	0.391229	0.527243	0.424889
0.578440	0.593747	0.641458	0.348784
0.595912	0.591881	0.433247	0.385875
0.568390	0.595302	0.243125	0.383931
0.525625	0.421310	0.518364	0.497079
0.536347	0.519604	0.496837	0.357837
0.567237	0.505327	0.378893	0.365750
0.516451	0.461785	0.280561	0.368968
0.535525	0.517521	0.490223	0.344180
0.548277	0.514908	0.109145	0.404535
0.536837	0.490723	0.483477	0.431994
0.552830	0.460916	0.542854	0.375604
0.596666	0.628196	0.523952	0.473126
0.619951	0.492341	0.462552	0.424473
0.524404	0.561009	0.360986	0.430441
0.543381	0.513132	0.508877	0.358517
0.609929	0.614706	0.217144	0.400274
0.540162	0.599211	0.582227	0.313021
0.551156	0.342648	0.426822	0.441985
0.519490	0.603000	0.500322	0.348195
0.584515	0.581989	0.197912	0.397236
0.506742	0.507226	0.718683	0.312467
0.575000	0.510948	0.412004	0.378656
0.562550	0.506473	0.505934	0.340014
0.567136	0.640978	0.286724	0.393550
0.573463	0.576815	0.365278	0.404420
0.500859	0.631011	0.380386	0.285880
0.591816	0.593793	0.491429	0.345156
0.571515	0.364627	0.585765	0.456314
0.528439	0.576724	0.400977	0.304197
0.565712	0.575847	0.450638	0.335614
0.551795	0.530373	0.216522	0.384768
0.572000	0.524522	0.379075	0.372487
0.542738	0.441303	0.460322	0.348510
0.586355	0.491397	0.302679	0.377799
0.544246	0.598518	0.281140	0.382757
0.620172	0.570979	0.384127	0.445120
0.588337	0.654627	0.239417	0.324289
0.575518	0.555545	0.659602	0.412833
0.533878	0.480957	0.441429	0.340319
0.633782	0.550665	0.261966	0.410399
0.646057	0.345871	0.396765	0.505200
0.600868	0.537695	0.599211	0.435831
0.618621	0.686463	0.398186	0.365586
0.583132	0.420352	0.637467	0.380627
0.509173	0.444438	0.615903	0.337977
0.585686	0.504639	0.509856	0.366821
0.589402	0.440032	0.279721	0.504505
0.650563	0.591478	0.619991	0.415295
0.517263	0.486308	0.562996	0.356558
0.549615	0.486650	0.736738	0.620539
0.486592	0.529161	0.659452	0.405366
0.622134	0.491205	0.639604	0.406336
0.571265	0.510720	0.536107	0.410159
0.625243	0.510115	0.369200	0.421666
0.576128	0.470506	0.448270	0.348276
0.520763	0.564302	0.370884	0.356413
0.639929	0.467515	0.579207	0.410603
0.581569	0.541550	0.326298	0.341968
0.561705	0.352955	0.214742	0.411725
0.568049	0.519738	0.180217	0.415384
0.499412	0.506819	0.498056	0.379931
0.593131	0.661366	0.297251	0.480453
0.488577	0.540339	0.618398	0.327922
0.557546	0.332663	0.497995	0.406344
0.552247	0.416661	0.320389	0.350327
0.564988	0.486747	0.449391	0.367602
0.505044	0.420180	0.270972	0.334494
0.610771	0.411661	0.251202	0.422653
0.560576	0.678105	0.465409	0.388791
0.581711	0.560163	0.312354	0.437526
0.600214	0.622986	0.526607	0.434461
0.574716	0.542095	0.616806	0.356831
0.587319	0.467595	0.565925	0.383531
0.583736	0.502642	0.237110	0.440597
0.532953	0.619386	0.537832	0.296423
0.548320	0.694212	0.563303	0.323727
0.573692	0.445113	0.463226	0.454336
0.520283	0.462231	0.432513	0.340841
0.626664	0.414999	0.745563	0.387560
0.489960	0.508598	0.475178	0.438257
0.596099	0.531519	0.404401	0.462850
0.595736	0.453837	0.352059	0.368473
0.609240	0.484174	0.557598	0.367286
0.432605	0.437355	0.466743	0.264925
0.610985	0.512786	0.151358	0.402562
0.551875	0.466964	0.407588	0.358845
0.590722	0.468212	0.546652	0.410199
0.524220	0.435545	0.361414	0.364959
0.574947	0.588340	0.216633	0.349461
0.627824	0.567842	0.597851	0.389081
0.523445	0.487777	0.378366	0.376605
0.546701	0.549048	0.448976	0.389472
0.555784	0.557621	0.575133	0.420817
0.611731	0.452633	0.736549	0.429878
0.572349	0.461915	0.494194	0.474881
0.494090	0.366941	0.166887	0.379249
0.594635	0.475703	0.416165	0.424432
0.516913	0.554506	0.456941	0.348317
0.506323	0.614308	0.511754	0.365003
0.608837	0.401671	0.662649	0.383282
0.624428	0.576252	0.242323	0.368772
0.493581	0.489407	0.336616	0.395375
0.637683	0.345094	0.343977	0.475863
0.557891	0.515493	0.362367	0.355014
0.600149	0.475806	0.362130	0.436949
0.614772	0.518369	0.260323	0.390381
0.530420	0.426987	0.593685	0.365131
0.586509	0.591584	0.453866	0.399472
0.486565	0.596888	0.386713	0.269330
0.593135	0.546580	0.297946	0.470051
0.568924	0.480317	0.568767	0.439368
0.607538	0.468002	0.218806	0.435260
0.557075	0.530728	0.275013	0.443548
0.534289	0.591090	0.605117	0.329683
0.602891	0.580409	0.606372	0.499741
0.602800	0.608830	0.471229	0.418574
0.549299	0.489330	0.746713	0.457398
0.562753	0.533600	0.430055	0.383796
0.561728	0.571630	0.630067	0.393630
0.547937	0.577995	0.454164	0.345335
0.548964	0.406277	0.599925	0.341608
0.573800	0.489200	0.219664	0.419983
0.565365	0.480804	0.312869	0.471591
0.537270	0.419078	0.309765	0.405331
0.552349	0.505737	0.422574	0.385080
0.570338	0.645489	0.512897	0.355823
0.582224	0.497307	0.342485	0.406508
0.585123	0.435252	0.537352	0.360977
0.501338	0.494974	0.494868	0.377366
0.612482	0.572990	0.335849	0.452217
0.611040	0.482659	0.496869	0.399082
0.593612	0.532425	0.369568	0.353265
0.549897	0.499741	0.494235	0.415699
0.553660	0.697663	0.275826	0.370401
0.519508	0.446756	0.551236	0.322601
0.534464	0.560232	0.561525	0.457813
0.588056	0.407286	0.238295	0.386648
0.491398	0.396001	0.375468	0.332373
0.538345	0.417919	0.271935	0.330854
0.535209	0.528152	0.577861	0.381198
0.533108	0.543121	0.564441	0.361355
0.599581	0.426920	0.546046	0.380079
0.490851	0.400809	0.514003	0.448213
0.490766	0.562125	0.480485	0.295870
0.541955	0.578145	0.539159	0.374193
0.559353	0.558057	0.509669	0.467666
0.544200	0.590686	0.324600	0.317828
0.585458	0.494953	0.550469	0.353813
0.530416	0.424768	0.447464	0.355099
0.628846	0.454791	0.763392	0.409491
0.571686	0.632332	0.301128	0.421015
0.490874	0.389448	0.269957	0.326642
0.597032	0.470846	0.488430	0.360596
0.584533	0.530301	0.538061	0.501153
0.643354	0.632040	0.406822	0.455190
0.510552	0.471465	0.332777	0.353729
0.561067	0.556847	0.268095	0.318533
0.553329	0.636164	0.558745	0.357411
0.569493	0.404097	0.236453	0.352751
0.547984	0.491583	0.450689	0.386638
0.495997	0.603132	0.438354	0.395250
0.547300	0.578062	0.486809	0.369810
0.499728	0.555465	0.706116	0.309242
0.564666	0.467109	0.307114	0.446097
0.508081	0.463114	0.470455	0.307105
0.575051	0.468098	0.719708	0.454120
0.490104	0.523473	0.504357	0.337835
0.497582	0.567142	0.342357	0.363289
0.568769	0.433209	0.266567	0.364073
0.575251	0.613702	0.697451	0.405556
0.651813	0.577696	0.449478	0.387901
0.577459	0.463328	0.543428	0.448756
0.490863	0.640102	0.590563	0.428993
0.624617	0.502524	0.474529	0.435977
0.626073	0.505874	0.431725	0.380728
0.527641	0.552841	0.481041	0.385298
0.528709	0.439293	0.455233	0.387441
0.564849	0.526071	0.268583	0.421776
0.528353	0.592400	0.381586	0.417179
0.584109	0.570213	0.641651	0.481478
0.618376	0.556653	0.303569	0.420672
0.523742	0.551104	0.359863	0.324726
0.526683	0.543941	0.540663	0.432171
0.533807	0.546650	0.504091	0.443599
0.538073	0.491449	0.464819	0.336245
0.617682	0.451507	0.671504	0.464895
0.512894	0.508128	0.534701	0.338421
0.583050	0.530061	0.639476	0.397791
0.525213	0.332942	0.546556	0.351366
0.624075	0.519160	0.399536	0.368530
0.564416	0.549603	0.458816	0.395234
0.567439	0.543872	0.519976	0.359248
0.594571	0.512430	0.404022	0.373244
0.591972	0.642796	0.370267	0.436718
0.574111	0.401299	0.494072	0.506438
0.589816	0.467251	0.554299	0.386687
0.515706	0.522710	0.547571	0.322878
0.515019	0.636986	0.615229	0.322980
0.535769	0.328875	0.241666	0.378564
0.540393	0.582325	0.444162	0.398538
0.590261	0.558209	0.427301	0.395713
0.574066	0.509182	0.614960	0.382659
0.599312	0.516797	0.671151	0.441323
0.588324	0.559518	0.481722	0.394191
0.589885	0.316704	0.438976	0.450873
0.618452	0.527558	0.341305	0.401275
0.542903	0.668116	0.599796	0.400072
0.517784	0.356873	0.629096	0.366386
0.579463	0.578589	0.584415	0.378314
0.560686	0.493167	0.601208	0.348839
0.521118	0.489961	0.353517	0.541164
0.586992	0.541231	0.349241	0.594398
0.555377	0.579670	0.302572	0.321856
0.606349	0.359019	0.645858	0.385120
0.582919	0.407904	0.347010	0.482633
0.562147	0.570591	0.519147	0.450273
0.513288	0.507069	0.399372	0.299717
0.593435	0.507464	0.266255	0.370804
0.585367	0.571670	0.537733	0.446984
0.577932	0.448550	0.289638	0.387725
0.581001	0.517518	0.323100	0.385280
0.533472	0.550338	0.432042	0.325665
0.538551	0.588601	0.517082	0.329411
0.660538	0.580122	0.733603	0.526262
0.532732	0.501438	0.355848	0.512565
0.588089	0.514608	0.409145	0.381671
0.515474	0.482619	0.383043	0.428639
0.618036	0.520337	0.466449	0.411973
0.533645	0.446967	0.305335	0.357105
0.563707	0.569710	0.545626	0.345739
0.603396	0.465455	0.592055	0.384604
0.599149	0.423497	0.442704	0.434588
0.562891	0.528719	0.666331	0.424731
0.493422	0.458125	0.445727	0.308536
0.579927	0.456141	0.459665	0.384936
0.498945	0.544885	0.348803	0.360193
0.587105	0.571351	0.432584	0.513585
0.490901	0.477767	0.602951	0.304871
0.529612	0.434799	0.390641	0.349944
0.607840	0.566110	0.456295	0.487024
0.508946	0.445314	0.257946	0.524299
0.511689	0.535618	0.706725	0.318617
0.564371	0.543873	0.451091	0.361299
0.600592	0.528706	0.296222	0.427848
0.502733	0.505443	0.590265	0.410091
0.598448	0.561326	0.496020	0.490025
0.484984	0.679005	0.294550	0.293374
0.537901	0.487922	0.389484	0.371262
0.599266	0.463409	0.542125	0.389814
0.561314	0.480554	0.558481	0.340764
0.566834	0.473601	0.452894	0.363901
0.543884	0.447236	0.328593	0.487985
0.527751	0.593003	0.390932	0.408637
0.620114	0.605999	0.520870	0.372430
0.626111	0.599294	0.317652	0.389138
0.596380	0.616795	0.591722	0.360791
0.597492	0.446476	0.543490	0.362613
0.549040	0.403394	0.423200	0.417689
0.555731	0.519441	0.514153	0.431963
0.606476	0.461520	0.486590	0.457693
0.610330	0.527829	0.174718	0.477844
0.597561	0.498602	0.266864	0.388993
0.551533	0.466013	0.558589	0.448777
0.568111	0.394434	0.559257	0.404390
0.531516	0.552877	0.173700	0.333629
0.540165	0.500094	0.355031	0.366955
0.559212	0.433665	0.215857	0.350223
0.617438	0.499045	0.308452	0.446021
0.471264	0.698079	0.358859	0.264354
0.565275	0.420899	0.765847	0.370419
0.640343	0.428643	0.562800	0.437793
0.593701	0.469208	0.275889	0.450056
0.583178	0.580357	0.610282	0.391479
0.631920	0.578126	0.134579	0.501790
0.541585	0.729807	0.418724	0.412705
0.527967	0.619335	0.577338	0.302856
0.579936	0.376640	0.294080	0.405448
0.598634	0.459125	0.475724	0.441901
0.483137	0.538000	0.365930	0.392536
0.565694	0.542025	0.520508	0.341692
0.526225	0.602883	0.212582	0.333371
0.507225	0.468131	0.395118	0.342098
0.580313	0.623910	0.309826	0.387768
0.606700	0.513213	0.450033	0.386419
0.526512	0.514964	0.362644	0.325683
0.553124	0.454533	0.352738	0.391041
0.496351	0.429370	0.243572	0.404269
0.588670	0.525608	0.494676	0.400917
0.602148	0.521631	0.262680	0.382780
0.519714	0.509485	0.405615	0.476276
0.560201	0.361612	0.401096	0.395626
0.605279	0.409255	0.445081	0.390239
0.515588	0.424018	0.613222	0.435870
0.581790	0.445559	0.327760	0.422207
0.563733	0.499686	0.605403	0.361704
0.596465	0.560619	0.514045	0.372105
0.577557	0.473267	0.563125	0.447225
0.517926	0.544825	0.584183	0.422015
0.501850	0.502416	0.578883	0.304487
0.534219	0.453101	0.555989	0.416597
0.505954	0.645913	0.436448	0.403422
0.559306	0.447705	0.732128	0.367004
0.591465	0.533821	0.339686	0.379350
0.604159	0.491927	0.580579	0.369236
0.535576	0.549537	0.319948	0.429729
0.497708	0.609746	0.389482	0.431068
0.547295	0.605867	0.309507	0.337583
0.495672	0.443868	0.693724	0.310847
0.576365	0.439234	0.296280	0.392973
0.511090	0.478061	0.105028	0.310484
0.581149	0.521291	0.385619	0.503625
0.576042	0.467438	0.682169	0.376400
0.587079	0.504873	0.383216	0.422352
0.521448	0.514712	0.363404	0.327423
0.588436	0.587838	0.469212	0.385960
0.568183	0.450531	0.280759	0.460239
0.587894	0.575438	0.365922	0.363227
0.521445	0.632112	0.698988	0.397325
0.558592	0.625575	0.460441	0.369895
0.628943	0.423898	0.430833	0.433557
0.568119	0.585642	0.267924	0.397045
0.575589	0.516404	0.610584	0.398182
0.569117	0.532096	0.630139	0.369330
0.526973	0.484421	0.308066	0.341486
0.593544	0.506993	0.503359	0.370292
0.545168	0.551836	0.426808	0.395195
0.569289	0.429892	0.560743	0.475632
0.519832	0.558945	0.487469	0.384259
0.472945	0.649546	0.489434	0.296086
0.550516	0.407563	0.757755	0.450901
0.537232	0.336470	0.286003	0.383918
0.549900	0.484906	0.428718	0.385593
0.550731	0.530395	0.447356	0.365574
0.647156	0.406382	0.567155	0.420163
0.561523	0.403589	0.622469	0.412063
0.535461	0.598155	0.516906	0.492193
0.584643	0.400065	0.285039	0.358638
0.579634	0.441891	0.416893	0.405457
0.562157	0.538831	0.087148	0.333729
0.607731	0.607886	0.595782	0.503814
0.449928	0.440485	0.275027	0.473266
0.595818	0.475725	0.421845	0.380615
0.486020	0.513961	0.301523	0.371567
0.533363	0.483522	0.280086	0.333939
0.630586	0.647702	0.487377	0.451239
0.573230	0.433595	0.418873	0.398858
0.573750	0.620890	0.422170	0.341460
0.526085	0.547224	0.730918	0.380343
0.598416	0.491436	0.381797	0.388996
0.553286	0.586953	0.657070	0.478730
0.536484	0.338970	0.339515	0.408024
0.482531	0.429934	0.438789	0.354578
0.560371	0.573521	0.219646	0.395326
0.577708	0.412281	0.639747	0.400856
0.479383	0.594091	0.397379	0.412915
0.555140	0.629773	0.287755	0.400102
0.615683	0.670491	0.693470	0.452214
0.524652	0.472220	0.544665	0.324342
0.632459	0.526488	0.215541	0.430973
0.622007	0.601875	0.358935	0.513185
0.518144	0.734469	0.459967	0.327763
0.575025	0.690791	0.526853	0.317688
0.550657	0.490120	0.365159	0.341264
0.495128	0.420478	0.279847	0.344709
0.528951	0.481303	0.516319	0.342591
0.492979	0.450235	0.543897	0.348870
0.622269	0.554148	0.168443	0.408213
0.628000	0.452938	0.482445	0.432162
0.590648	0.535519	0.167402	0.393948
0.565505	0.590306	0.500467	0.343421
0.570662	0.514893	0.311477	0.333358
0.564839	0.599876	0.458406	0.503383
0.594948	0.598472	0.565629	0.340719
0.577220	0.538446	0.443544	0.382395
0.510122	0.533652	0.236570	0.322759
0.587571	0.565939	0.668394	0.423611
0.581580	0.590961	0.625999	0.379332
0.541913	0.529786	0.359740	0.361381
0.567782	0.387471	0.147896	0.478678
0.617233	0.570723	0.449280	0.357552
0.508690	0.530353	0.418715	0.293553
0.602074	0.639142	0.546897	0.387420
0.528577	0.366744	0.557153	0.434246
0.598608	0.554389	0.418867	0.417546
0.546664	0.456526	0.476466	0.385290
0.585387	0.589533	0.514514	0.349059
0.547813	0.393222	0.312438	0.371700
0.582455	0.518407	0.276209	0.400709
0.542349	0.560656	0.219663	0.557972
0.569191	0.501281	0.567943	0.379657
0.527569	0.542406	0.683700	0.358329
0.593051	0.637403	0.328077	0.336928
0.578142	0.534052	0.437775	0.363246
0.527365	0.465604	0.543121	0.434452
0.567396	0.594611	0.550338	0.365455
0.511618	0.473710	0.396562	0.330269
0.612377	0.488238	0.714837	0.410221
0.555084	0.465642	0.563058	0.404749
0.609896	0.636431	0.654579	0.615310
0.606337	0.548339	0.565949	0.495951
0.618120	0.657428	0.398771	0.454908
0.553393	0.513717	0.364810	0.325718
0.596607	0.444858	0.174574	0.434681
0.490702	0.528761	0.410482	0.369817
0.559278	0.465793	0.298727	0.358194
0.607246	0.437035	0.462514	0.457969
0.613361	0.447530	0.534498	0.500658
0.575197	0.553538	0.494747	0.352937
0.506982	0.558702	0.574444	0.337352
0.573772	0.650519	0.647364	0.430853
0.446771	0.468792	0.403703	0.325985
0.682064	0.430873	0.560844	0.525355
0.572047	0.508009	0.410942	0.473610
0.595141	0.433518	0.332475	0.429671
0.606942	0.517148	0.791387	0.435231
0.560442	0.553116	0.397285	0.402392
0.544562	0.419593	0.502749	0.356990
0.597125	0.561554	0.576122	0.424094
0.490027	0.435568	0.555517	0.346956
0.546952	0.510416	0.443524	0.336265
0.591791	0.593710	0.501485	0.459667
0.532868	0.488059	0.366681	0.328216
0.546307	0.525258	0.427662	0.378000
0.533887	0.441756	0.525259	0.363430
0.607622	0.465263	0.254740	0.375347
0.591627	0.548863	0.461039	0.464351
0.535649	0.554080	0.673486	0.357191
0.551744	0.490316	0.460771	0.488050
0.595160	0.451768	0.355959	0.369678
0.563841	0.430388	0.481973	0.390029
0.570477	0.506897	0.500169	0.347958
0.603150	0.489298	0.289100	0.408043
0.647829	0.419403	0.481845	0.494276
0.354064	0.544199	0.441257	0.254507
0.629351	0.577569	0.452330	0.339388
0.741001	0.706396	0.462884	0.483887
0.751944	0.773470	0.419032	0.516694
0.641252	0.496715	0.456512	0.556208
0.782716	0.499538	0.445970	0.391451
0.784753	0.341168	0.476957	0.268222
0.535035	0.548210	0.409158	0.398885
0.658566	0.361118	0.351917	0.500822
0.580986	0.494724	0.452799	0.402581
0.415690	0.707608	0.496883	0.358319
0.550675	0.461727	0.482491	0.256571
0.443808	0.299959	0.460931	0.378269
0.612915	0.327353	0.351250	0.489529
0.383987	0.400592	0.439381	0.352860
0.854988	0.533630	0.452692	0.541186
0.407188	0.462891	0.483435	0.121341
0.611759	0.431982	0.438477	0.429946
0.663276	0.542058	0.458229	0.440395
0.571262	0.459890	0.395416	0.516509
0.320005	0.523469	0.412007	0.300947
0.740557	0.584985	0.458930	0.156142
0.749286	0.449663	0.502440	0.435050
0.573191	0.574344	0.393147	0.417986
0.429367	0.687188	0.381019	0.295816
0.603360	0.524885	0.378022	0.380140
0.453907	0.572974	0.458320	0.436512
0.673245	0.591167	0.450605	0.527902
0.625888	0.357305	0.423621	0.370617
0.454697	0.466931	0.480547	0.448676
0.590779	0.505710	0.507012	0.442921
0.524816	0.714081	0.360696	0.340586
0.236557	0.575674	0.409481	0.243260
0.502055	0.430983	0.366474	0.488242
0.707043	0.695447	0.374669	0.537921
0.440979	0.463121	0.412339	0.449549
0.472028	0.510001	0.437182	0.353652
0.520841	0.356091	0.504279	0.315255
0.409950	0.463992	0.443312	0.399105
0.438870	0.554385	0.430044	0.164881
0.564752	0.572325	0.395261	0.407837
0.533647	0.624859	0.398468	0.342660
0.638427	0.613344	0.383521	0.454675
0.611991	0.557241	0.372310	0.253331
0.794991	0.553589	0.424676	0.425870
0.729089	0.696582	0.528260	0.360950
0.676716	0.616881	0.440067	0.251811
0.696763	0.439566	0.540173	0.416471
0.470635	0.582424	0.372923	0.307699
0.620216	0.672798	0.372616	0.522598
0.317305	0.639044	0.390823	0.328197
0.666992	0.406049	0.394038	0.567698
0.394827	0.407145	0.426078	0.432237
0.482715	0.726321	0.462740	0.374122
0.407801	0.629546	0.450890	0.277058
0.758765	0.665033	0.461235	0.551953
0.684766	0.269900	0.503828	0.346612
0.525270	0.500185	0.428943	0.246335
0.582039	0.343275	0.364546	0.395815
0.602480	0.255887	0.417236	0.322594
0.616216	0.469198	0.520460	0.417445
0.354859	0.561781	0.462774	0.302158
0.734343	0.550777	0.486159	0.408879
0.397324	0.591377	0.424453	0.359174
0.486651	0.607973	0.437246	0.435456
0.526060	0.405089	0.323380	0.418630
0.585217	0.440928	0.483302	0.471171
0.502975	0.465917	0.479132	0.325249
0.501391	0.753167	0.427555	0.304615
0.492540	0.729554	0.485876	0.373102
0.598419	0.447784	0.353633	0.467876
0.359571	0.534145	0.485826	0.323812
0.694621	0.248050	0.440479	0.568745
0.473622	0.346675	0.473975	0.482427
0.565985	0.734677	0.477327	0.471927
0.450575	0.574736	0.480449	0.304980
0.607677	0.572954	0.441434	0.274340
0.549336	0.560606	0.568327	0.477486
0.589339	0.486977	0.395368	0.498923
0.645224	0.646235	0.444184	0.413394
0.435400	0.520493	0.487927	0.172782
0.453388	0.577636	0.411880	0.421792
0.579776	0.691043	0.448016	0.405807
0.474691	0.635053	0.360203	0.361830
0.354369	0.543109	0.401982	0.364519
0.416931	0.320323	0.394185	0.391627
0.569133	0.517494	0.355225	0.475831
0.595497	0.492477	0.435186	0.460765
0.632641	0.503919	0.450301	0.472679
0.469919	0.424382	0.389905	0.360866
0.590264	0.495694	0.426407	0.377108
0.491298	0.474665	0.380793	0.338805
0.445194	0.177777	0.452900	0.434508
0.568592	0.494337	0.476230	0.522241
0.724512	0.347147	0.518812	0.313103
0.497482	0.449962	0.442397	0.344566
0.325721	0.298400	0.499059	0.388386
0.407204	0.523178	0.425461	0.337000
0.697879	0.361162	0.509132	0.460582
0.429872	0.410247	0.389484	0.362369
0.631734	0.724538	0.419902	0.410026
0.330724	0.603018	0.376077	0.341874
0.392230	0.357496	0.392175	0.402602
0.582400	0.421343	0.479025	0.406632
0.599619	0.414280	0.480806	0.257467
0.654734	0.556396	0.438389	0.505373
0.757858	0.316764	0.342006	0.569336
0.688587	0.330806	0.407080	0.361278
0.318972	0.366258	0.471806	0.291541
0.694369	0.560075	0.382332	0.484656
0.496931	0.468501	0.376181	0.326297
0.553696	0.691310	0.419106	0.463659
0.510240	0.525628	0.480507	0.318634
0.611778	0.451130	0.431043	0.452224
0.601386	0.626205	0.525829	0.376049
0.898040	0.577991	0.532395	0.624026
0.483168	0.428504	0.411995	0.386837
0.574948	0.404100	0.418567	0.194405
0.568960	0.336135	0.506231	0.474703
0.660223	0.522911	0.426283	0.373887
0.906032	0.562367	0.381214	0.435961
0.624491	0.473808	0.484624	0.396484
0.448138	0.524764	0.305470	0.421171
0.694135	0.471929	0.508365	0.464644
0.571692	0.534669	0.429068	0.446824
0.544149	0.309829	0.421836	0.399253
0.632259	0.559293	0.496066	0.480355
0.517313	0.531505	0.457442	0.463094
0.664887	0.247064	0.495473	0.588205
0.429085	0.651433	0.451248	0.249042
0.701614	0.326158	0.395398	0.394970
0.637959	0.513277	0.412490	0.404457
0.623391	0.474535	0.449422	0.520418
0.462019	0.515139	0.523980	0.428895
0.537217	0.650610	0.430233	0.427065
0.630857	0.478115	0.428856	0.301176
0.595254	0.706333	0.461822	0.466662
0.772060	0.408798	0.528128	0.603781
0.581773	0.427800	0.425316	0.408029
0.213645	0.597749	0.441557	0.257160
0.872544	0.435155	0.423716	0.670146
0.309397	0.674235	0.435044	0.289569
0.515211	0.431178	0.522077	0.422531
0.414339	0.501684	0.435237	0.319572
0.516782	0.526532	0.442297	0.383817
0.603863	0.513421	0.484738	0.428541
0.534918	0.602117	0.468516	0.351887
0.655014	0.496123	0.470616	0.557140
0.841536	0.533963	0.486329	0.407277
0.651202	0.549454	0.406212	0.447183
0.266987	0.881498	0.454945	0.273260
0.705974	0.458396	0.471509	0.390242
0.567852	0.488866	0.484861	0.418032
0.618276	0.710871	0.493805	0.452111
0.479162	0.528548	0.465425	0.255005
0.727191	0.385694	0.493946	0.375321
0.595419	0.313353	0.435796	0.512959
0.465868	0.521375	0.512726	0.454911
0.517697	0.291986	0.407867	0.313550
0.570164	0.487276	0.454413	0.492478
0.676121	0.445513	0.395104	0.436691
0.524673	0.432964	0.442610	0.438555
0.557246	0.342907	0.427594	0.365535
0.465536	0.791737	0.504431	0.210475
0.843516	0.481387	0.458277	0.339324
0.404810	0.686539	0.415464	0.316923
0.753612	0.392503	0.481983	0.317383
0.665624	0.675177	0.414907	0.482024
0.655303	0.543475	0.416318	0.415417
0.455555	0.387710	0.360047	0.238502
0.488130	0.482774	0.444607	0.451558
0.490477	0.455799	0.432239	0.468902
0.791565	0.296261	0.392795	0.409915
0.560810	0.545636	0.515496	0.330781
0.261234	0.454926	0.442574	0.267025
0.458733	0.727806	0.500452	0.368217
0.545976	0.419584	0.398730	0.414986
0.354671	0.598079	0.421160	0.288178
0.557069	0.502064	0.462496	0.357298
0.697960	0.453862	0.435607	0.464301
0.424757	0.739733	0.482493	0.359329
0.787778	0.436223	0.411038	0.355527
0.454709	0.547634	0.502888	0.433988
0.684337	0.529032	0.443349	0.521762
0.441613	0.512462	0.523565	0.324889
0.580143	0.354904	0.386839	0.266843
0.605029	0.550135	0.525087	0.427620
0.450038	0.557322	0.487536	0.379604
0.504020	0.498881	0.486630	0.405400
0.452465	0.349640	0.432293	0.413287
0.735952	0.581304	0.480068	0.417389
0.560557	0.434808	0.525573	0.519182
0.651297	0.560085	0.484778	0.547689
0.552279	0.521309	0.489370	0.336634
0.351090	0.451244	0.443974	0.208644
0.541689	0.415569	0.485460	0.416467
0.344941	0.497561	0.438232	0.205542
0.817636	0.460256	0.451672	0.372134
0.457341	0.537823	0.495519	0.378316
0.536368	0.371532	0.481892	0.449296
0.621543	0.390625	0.489991	0.492051
0.580372	0.532773	0.453365	0.451227
0.533746	0.435328	0.437907	0.400422
0.566691	0.723772	0.432612	0.359343
0.405952	0.745432	0.483624	0.326874
0.728765	0.550639	0.375560	0.537609
0.502324	0.299735	0.478857	0.437189
0.340517	0.504285	0.467926	0.366522
0.540887	0.619296	0.438933	0.336711
0.607325	0.636868	0.413408	0.205624
0.532567	0.483849	0.404689	0.331147
0.649498	0.231260	0.386574	0.435677
0.505391	0.465479	0.399475	0.402084
0.696754	0.481083	0.497157	0.465602
0.612276	0.543958	0.499999	0.332286
0.712513	0.459854	0.437555	0.565222
0.539562	0.613353	0.443413	0.419933
0.609571	0.602372	0.351607	0.494354
0.368771	0.541358	0.524642	0.300574
0.439013	0.694463	0.383758	0.191097
0.464272	0.595599	0.371441	0.362690
0.527998	0.527759	0.409873	0.421444
0.620263	0.491200	0.435258	0.484025
0.774702	0.572135	0.449154	0.490287
0.752082	0.493981	0.488263	0.438150
0.842387	0.664856	0.447985	0.232159
0.401395	0.460638	0.481363	0.241230
0.387708	0.560831	0.437954	0.355364
0.377069	0.601237	0.410265	0.354197
0.489667	0.568296	0.422757	0.312463
0.566981	0.618141	0.495993	0.348404
0.443743	0.627738	0.395615	0.317158
0.454154	0.388852	0.412873	0.364189
0.688895	0.597625	0.491157	0.526144
0.748909	0.502235	0.464967	0.457748
0.645128	0.674855	0.488500	0.392102
0.644644	0.348121	0.530498	0.436287
0.643094	0.582486	0.455742	0.332682
0.716009	0.326296	0.435530	0.637667
0.470275	0.429509	0.477255	0.284266
0.391890	0.324623	0.449757	0.270546
0.505108	0.434639	0.464030	0.342113
0.597590	0.742139	0.439864	0.223896
0.398690	0.544240	0.531194	0.276550
0.429423	0.468563	0.498178	0.367019
0.362121	0.575664	0.497255	0.150790
0.426202	0.776244	0.483561	0.386262
0.807268	0.678072	0.454645	0.610139
0.575304	0.339430	0.443011	0.458612
0.760161	0.466343	0.543894	0.431041
0.411310	0.773850	0.443441	0.334620
0.383435	0.509199	0.480705	0.373439
0.568306	0.577556	0.474459	0.411902
0.546522	0.369226	0.395845	0.455658
0.818692	0.519590	0.481528	0.292542
0.718305	0.524440	0.427770	0.535171
0.511200	0.539316	0.370674	0.464091
0.544152	0.498848	0.462498	0.428146
0.693832	0.620985	0.461894	0.517637
0.297647	0.518416	0.464902	0.206191
0.764777	0.559472	0.502071	0.569511
0.647471	0.481480	0.489512	0.346469
0.502537	0.571926	0.517691	0.398192
0.417917	0.687369	0.411808	0.223083
0.688588	0.574100	0.457129	0.400707
0.620293	0.444036	0.449776	0.346235
0.481341	0.352433	0.426075	0.471095
0.563689	0.504081	0.448081	0.517187
0.500025	0.503051	0.344099	0.428304
0.566589	0.673040	0.431284	0.323946
0.908805	0.542974	0.597634	0.275158
0.529689	0.613105	0.449963	0.383506
0.506285	0.498360	0.400012	0.333696
0.320164	0.463368	0.459381	0.370307
0.498730	0.484414	0.565503	0.395128
0.557631	0.567961	0.430374	0.418318
0.401530	0.358977	0.448252	0.428414
0.597417	0.529227	0.444741	0.401719
0.550217	0.448604	0.409854	0.473153
0.424284	0.502062	0.447421	0.416975
0.541916	0.302462	0.371920	0.489449
0.614901	0.647099	0.426393	0.273656
0.566029	0.317818	0.490201	0.488514
0.529546	0.517064	0.436677	0.445653
0.457955	0.651197	0.456934	0.357449
0.685451	0.290096	0.376996	0.456339
0.468564	0.526156	0.414405	0.282654
0.673716	0.402882	0.360967	0.493961
0.555960	0.432866	0.395797	0.512231
0.540635	0.717054	0.356895	0.263288
0.607156	0.604223	0.422916	0.438311
0.372689	0.238134	0.399517	0.312899
0.450745	0.427143	0.424987	0.369510
0.585371	0.322455	0.382376	0.495459
0.563725	0.612754	0.437340	0.377591
0.511083	0.537427	0.433872	0.400486
0.372659	0.306341	0.477677	0.353264
0.525744	0.540819	0.410825	0.238929
0.469664	0.556721	0.579059	0.376587
0.683888	0.461155	0.453635	0.498044
0.595232	0.555513	0.473289	0.467886
0.640704	0.593448	0.391636	0.478846
0.596986	0.571637	0.373486	0.261033
0.411046	0.633390	0.447230	0.378967
0.546131	0.498933	0.464253	0.426150
0.459217	0.518469	0.430900	0.337391
0.503640	0.463343	0.443411	0.486200
0.674853	0.401301	0.474490	0.413592
0.499866	0.549169	0.460839	0.449449
0.667666	0.565609	0.437320	0.539138
0.571761	0.477958	0.469104	0.523949
0.691920	0.815029	0.429256	0.534227
0.505450	0.434831	0.444605	0.321310
0.438944	0.585979	0.469991	0.418699
0.394967	0.417833	0.490596	0.305238
0.754863	0.518934	0.474413	0.470419
0.458882	0.616000	0.448399	0.375368
0.431331	0.511447	0.442266	0.319382
0.552755	0.582639	0.355132	0.286965
0.531787	0.479362	0.459945	0.409069
0.592913	0.553729	0.478795	0.274202
0.532549	0.516002	0.497337	0.323815
0.586746	0.572526	0.471500	0.388328
0.647374	0.453153	0.447985	0.394504
0.415078	0.509294	0.395143	0.311389
0.563877	0.554340	0.494883	0.367660
0.616595	0.492323	0.385544	0.242440
0.457738	0.581160	0.420736	0.358491
0.580707	0.675485	0.494668	0.403273
0.703650	0.262407	0.414582	0.384367
0.731822	0.519833	0.465964	0.557528
0.538124	0.821601	0.443423	0.139226
0.714479	0.666986	0.508035	0.558065
0.645413	0.432760	0.473511	0.406688
0.462150	0.573192	0.502480	0.439003
0.761314	0.564571	0.403263	0.527916
0.407770	0.436978	0.460221	0.411311
0.732990	0.594176	0.464492	0.548174
0.389378	0.672509	0.361805	0.355181
0.287287	0.310239	0.435614	0.327725
0.360205	0.622287	0.381995	0.357942
0.495689	0.552841	0.457510	0.396554
0.759666	0.462056	0.395899	0.425121
0.276391	0.474840	0.400025	0.266054
0.467663	0.573832	0.469531	0.447235
0.397063	0.430503	0.425990	0.396822
0.516403	0.437703	0.462721	0.471167
0.482204	0.446962	0.406592	0.378074
0.507531	0.511717	0.510150	0.371045
0.667548	0.716392	0.448003	0.401891
0.605978	0.503210	0.399910	0.175146
0.442156	0.679203	0.382588	0.090334
0.472924	0.438372	0.448474	0.373852
0.653479	0.502393	0.438601	0.369944
0.717561	0.397248	0.517604	0.379708
0.556963	0.447222	0.355099	0.493867
0.578626	0.474801	0.472314	0.434876
0.535005	0.277412	0.530719	0.468179
0.621391	0.235377	0.507244	0.529173
0.549668	0.471801	0.517827	0.418747
0.358538	0.579232	0.393679	0.307801
0.538353	0.576467	0.505279	0.489497
0.690872	0.559454	0.500132	0.480649
0.474484	0.375913	0.437079	0.364573
0.665554	0.529812	0.484775	0.424389
0.545120	0.239368	0.429382	0.328717
0.342229	0.539864	0.332095	0.232431
0.601234	0.468768	0.377141	0.292166
0.381117	0.572116	0.450453	0.332318
0.739867	0.452514	0.493392	0.378226
0.453226	0.783711	0.437121	0.373937
0.506579	0.503424	0.382616	0.160234
0.603910	0.449448	0.461658	0.423276
0.417438	0.466593	0.477118	0.413765
0.447169	0.571166	0.444960	0.350727
0.438950	0.574969	0.497876	0.269854
0.631174	0.727056	0.491124	0.391504
0.553465	0.336634	0.405763	0.159371
0.469521	0.542119	0.424142	0.436242
0.527004	0.561169	0.439173	0.376457
0.412190	0.586441	0.422421	0.376717
0.547822	0.608266	0.406202	0.355530
0.340417	0.497391	0.442936	0.326161
0.617394	0.513243	0.493796	0.476810
0.435655	0.453949	0.447878	0.370949
0.521196	0.577376	0.434048	0.402790
0.861377	0.572723	0.522868	0.426059
0.754803	0.545833	0.458642	0.363124
0.694815	0.478366	0.521020	0.313612
0.604466	0.591983	0.460805	0.471287
0.510326	0.390780	0.472541	0.470663
0.671300	0.595195	0.389252	0.487977
0.696678	0.461756	0.421118	0.569570
0.550821	0.553331	0.378741	0.372617
0.632017	0.730603	0.436421	0.336514
0.589059	0.313307	0.399912	0.377809
0.529457	0.439530	0.439539	0.354875
0.596435	0.483042	0.441332	0.428352
0.534848	0.475885	0.490129	0.094087
0.642360	0.409521	0.437582	0.572571
0.543735	0.514115	0.408883	0.233865
0.574349	0.526795	0.449028	0.300917
0.431887	0.579832	0.449577	0.342038
0.628165	0.470436	0.476321	0.479383
0.593703	0.452856	0.412558	0.404502
0.467946	0.455973	0.424397	0.290858
0.867583	0.504304	0.400998	0.329276
0.542402	0.564994	0.439257	0.360567
0.586185	0.477144	0.471833	0.417012
0.628883	0.510452	0.335216	0.528232
0.561856	0.639913	0.408121	0.476904
0.766691	0.524139	0.456782	0.439480
0.457021	0.557178	0.401989	0.395590
0.494943	0.605103	0.474215	0.324252
0.513238	0.615530	0.476915	0.468404
0.505719	0.475992	0.482243	0.360725
0.757582	0.445925	0.392012	0.464807
0.597668	0.508405	0.387421	0.253702
0.710098	0.439233	0.444348	0.214327
0.798215	0.424848	0.572947	0.479312
0.446928	0.678443	0.499438	0.381596
0.585959	0.507911	0.377035	0.351546
0.599553	0.521497	0.490939	0.344198
0.450896	0.558644	0.433104	0.432599
0.506860	0.523121	0.478242	0.287662
0.425916	0.555801	0.465108	0.315147
0.970445	0.244693	0.394554	0.517786
0.681414	0.264341	0.474787	0.468596
0.502169	0.175293	0.444562	0.442673
0.664671	0.438058	0.411105	0.577969
0.621589	0.676815	0.396741	0.338790
0.494504	0.611139	0.465694	0.423779
0.358587	0.281209	0.428377	0.426630
0.375551	0.522834	0.441591	0.323807
0.815647	0.374245	0.394741	0.636603
0.169991	0.452028	0.551227	0.175301
0.547752	0.457048	0.477201	0.417450
0.596239	0.643514	0.365267	0.394764
0.537699	0.516336	0.450818	0.056056
0.644141	0.693230	0.469771	0.445927
0.618177	0.501498	0.450055	0.441965
0.644976	0.408164	0.439145	0.547387
0.567876	0.481625	0.369626	0.298584
0.464595	0.410341	0.463126	0.447410
0.505721	0.461094	0.435145	0.402045
0.665554	0.552667	0.412563	0.442632
0.685672	0.524098	0.448408	0.572245
0.555116	0.496138	0.424945	0.484883
0.643069	0.333545	0.406070	0.450937
0.536268	0.521144	0.426477	0.424458
0.642429	0.372969	0.468972	0.369287
0.560924	0.139797	0.459624	0.555818
0.527142	0.576358	0.466205	0.428601
0.677593	0.370348	0.431325	0.284378
0.512408	0.355024	0.433499	0.424921
0.361232	0.568667	0.410186	0.372212
0.714554	0.593718	0.382646	0.501263
0.690768	0.567822	0.463959	0.493243
0.340812	0.599226	0.436809	0.368338
0.580678	0.359960	0.400934	0.352775
0.463470	0.468630	0.475714	0.220043
0.409566	0.703892	0.420363	0.211166
0.699045	0.580030	0.468398	0.394822
0.583948	0.564567	0.456713	0.402392
0.598272	0.352416	0.432459	0.441322
0.469852	0.546811	0.463531	0.223813
0.661514	0.465408	0.400957	0.512221
0.376251	0.615774	0.516980	0.198266
0.710145	0.406085	0.481889	0.354335
0.299090	0.296441	0.445048	0.254041
0.764292	0.739441	0.415975	0.500164
0.412234	0.463591	0.434891	0.311002
0.670166	0.575779	0.464387	0.494643
0.682837	0.508672	0.434440	0.431540
0.383983	0.370828	0.456644	0.313244
0.619425	0.462077	0.418967	0.368572
0.598832	0.334295	0.369450	0.545482
0.745579	0.522311	0.467110	0.589590
0.819910	0.509510	0.440894	0.304615
0.562493	0.334639	0.502271	0.331870
0.441013	0.686738	0.436795	0.390068
0.457524	0.624492	0.472324	0.293638
0.402408	0.350662	0.401367	0.436126
0.642727	0.491181	0.486134	0.423979
0.574952	0.436741	0.481335	0.535709
0.520304	0.536007	0.393278	0.421510
0.922563	0.662989	0.451512	0.653959
0.547855	0.670878	0.411618	0.364980
0.528126	0.470479	0.402930	0.383439
0.641314	0.434253	0.454447	0.484892
0.609567	0.579893	0.528379	0.453235
0.465809	0.320769	0.347875	0.269252
0.509123	0.514301	0.442844	0.267842
0.218358	0.534064	0.504491	0.248405
0.435072	0.648857	0.461072	0.412082
0.692313	0.268443	0.500794	0.395402
0.395925	0.453320	0.489854	0.103936
0.533784	0.660077	0.417942	0.370707
0.652472	0.463839	0.437060	0.493973
0.583753	0.400152	0.425102	0.328050
0.552502	0.327179	0.373998	0.504513
0.651733	0.422482	0.446449	0.340914
0.658831	0.503927	0.539225	0.456198
0.405276	0.430493	0.508339	0.250157
0.777437	0.522454	0.385987	0.246470
0.610961	0.619936	0.473057	0.381970
0.661283	0.374728	0.395013	0.299358
0.470971	0.691609	0.509753	0.271446
0.477812	0.431114	0.499006	0.466016
0.681231	0.520888	0.477399	0.587118
0.637065	0.449735	0.423786	0.333217
0.283865	0.436116	0.314005	0.135909
0.593880	0.511887	0.418708	0.488367
0.640108	0.875524	0.388726	0.460717
0.547336	0.300078	0.414210	0.531986
0.503231	0.435206	0.373431	0.383486
0.489461	0.441436	0.456828	0.412721
0.326404	0.320345	0.505645	0.330070
0.438648	0.660768	0.375998	0.325131
0.409192	0.511967	0.356527	0.385132
0.318627	0.470681	0.490419	0.306589
0.506562	0.530046	0.370761	0.455683
0.509237	0.588961	0.463030	0.388310
0.715128	0.378965	0.490307	0.620173
0.354867	0.561727	0.389406	0.358217
0.320694	0.546190	0.484836	0.236658
0.494571	0.604162	0.447287	0.458877
0.426965	0.557627	0.472812	0.394437
0.589326	0.505716	0.545529	0.402920
0.464251	0.396442	0.437186	0.343162
0.651209	0.629901	0.471979	0.435614
0.637535	0.483152	0.416100	0.546245
0.375323	0.329017	0.404910	0.254697
0.659150	0.292325	0.528056	0.299856
0.672006	0.417499	0.445695	0.380879
0.414392	0.663269	0.378790	0.107288
0.398733	0.532709	0.484729	0.402371
0.437942	0.481697	0.450147	0.322477
0.420058	0.398334	0.602445	0.430854
1.000000	0.552094	0.491996	0.492282
0.781148	0.513618	0.510812	0.429541
0.669493	0.500586	0.459446	0.415198
0.415417	0.461061	0.505024	0.352302
0.608162	0.357295	0.418702	0.476591
0.733831	0.609558	0.475322	0.557098
0.565294	0.544164	0.409915	0.370226
0.753220	0.670460	0.436861	0.561099
0.257017	0.399185	0.443502	0.319195
0.543915	0.485421	0.458032	0.405441
0.772830	0.288643	0.457882	0.475111
0.438734	0.548154	0.404866	0.418997
0.747815	0.607569	0.427575	0.452640
0.634231	0.446015	0.424668	0.418058
0.580907	0.415761	0.368674	0.529825
0.331935	0.327256	0.425405	0.384846
0.369686	0.473521	0.509781	0.334685
0.707043	0.625113	0.486250	0.262798
0.511839	0.353408	0.547069	0.340441
0.599810	0.611715	0.446700	0.373221
0.391351	0.653466	0.442636	0.367694
0.566195	0.653910	0.424171	0.311134
0.574420	0.401863	0.475449	0.532009
0.507829	0.534427	0.444905	0.272530
0.699683	0.536197	0.526487	0.356662
0.570883	0.370947	0.530372	0.462452
0.676953	0.724067	0.469241	0.268437
0.587703	0.242111	0.421889	0.461093
0.383703	0.590504	0.472956	0.236628
0.640442	0.608618	0.406891	0.367128
0.783867	0.440705	0.479564	0.649454
0.522177	0.623177	0.417176	0.438581
0.764484	0.569524	0.462135	0.425189
0.684134	0.533922	0.493814	0.481451
0.549006	0.693790	0.504168	0.352260
0.552627	0.651126	0.429918	0.393738
0.334497	0.512483	0.436177	0.324247
0.603274	0.695668	0.446062	0.460435
0.479345	0.701374	0.428747	0.364833
0.432575	0.401769	0.500924	0.418273
0.824989	0.392739	0.367088	0.276818
0.518999	0.272808	0.408797	0.311723
0.462817	0.332689	0.479792	0.322392
0.826115	0.362319	0.433363	0.562878
0.406008	0.417656	0.381266	0.348051
0.501404	0.657960	0.424770	0.265136
0.619647	0.476260	0.442347	0.354298
0.414970	0.452763	0.454056	0.245114
0.756313	0.498692	0.451258	0.261276
0.507714	0.533812	0.415593	0.375291
0.859916	0.822823	0.434719	0.303367
0.541856	0.735922	0.468309	0.430848
0.606855	0.527479	0.452283	0.468607
0.518265	0.606290	0.431182	0.340404
0.413304	0.439698	0.508718	0.404649
0.357332	0.576891	0.386821	0.329584
0.794282	0.696074	0.458523	0.365951
0.926504	0.425588	0.426411	0.370266
0.543114	0.361569	0.421807	0.525408
0.500013	0.403328	0.386660	0.337135
0.516404	0.435893	0.420466	0.446913
0.595327	0.712100	0.443876	0.487733
0.452154	0.320793	0.465113	0.473906
0.509257	0.255219	0.449160	0.304509
0.822478	0.432036	0.476209	0.293629
0.603073	0.569152	0.512709	0.481989
0.321248	0.673326	0.432729	0.343299
0.415850	0.510681	0.352542	0.341485
0.618267	0.365229	0.481628	0.269863
0.443296	0.474205	0.424647	0.258488
0.632510	0.627089	0.481863	0.399868
0.440091	0.340359	0.317200	0.380861
0.505061	0.616828	0.484082	0.462243
0.427678	0.527629	0.416652	0.308997
0.689847	0.518810	0.433574	0.332466
0.516612	0.355202	0.461443	0.215988
0.668385	0.394182	0.484823	0.416677
0.592185	0.500639	0.412588	0.472904
0.549928	0.339009	0.410991	0.298798
0.383155	0.623705	0.478421	0.338876
0.710510	0.621755	0.413817	0.475272
0.409327	0.521435	0.419310	0.404439
0.592651	0.469959	0.482067	0.368339
0.621577	0.333738	0.388177	0.497411
0.578818	0.474522	0.357938	0.499968
0.556400	0.333807	0.389699	0.509733
0.624482	0.726069	0.535506	0.437935
0.403462	0.808250	0.486235	0.362389
0.470142	0.508129	0.469622	0.455048
0.481899	0.367940	0.516871	0.489770
0.700169	0.318556	0.455542	0.501785
0.372400	0.576408	0.431975	0.299574
0.577827	0.605409	0.432708	0.323250
0.555120	0.512773	0.463886	0.442430
0.629832	0.566740	0.430825	0.450752
0.599884	0.411254	0.366017	0.339559
0.528892	0.525246	0.462555	0.458061
0.521968	0.487267	0.417528	0.453283
0.447509	0.481016	0.365810	0.411278
0.402561	0.379372	0.482685	0.412377
0.362141	0.329922	0.434656	0.340915
0.654024	0.581930	0.432670	0.495037
0.745046	0.295649	0.512770	0.456662
0.582753	0.605041	0.403421	0.422581
0.527260	0.353408	0.533310	0.275718
0.473416	0.424346	0.475562	0.415372
0.506903	0.699462	0.487540	0.405691
0.537236	0.477186	0.423791	0.391087
0.520974	0.391155	0.473340	0.436168
0.597111	0.422836	0.478256	0.532311
0.661213	0.432411	0.499820	0.578287
0.564724	0.634124	0.462109	0.493073
0.617906	0.721089	0.448707	0.348369
0.713875	0.538334	0.485431	0.458502
0.500247	0.628303	0.533451	0.389177
0.411406	0.384522	0.357745	0.270198
0.706781	0.530882	0.376300	0.379081
0.425315	0.494678	0.383918	0.382169
0.635607	0.501629	0.382126	0.520425
0.572941	0.440572	0.406464	0.440753
0.703133	0.493316	0.425955	0.477198
0.551998	0.360325	0.467078	0.175542
0.527216	0.574535	0.342998	0.424507
0.270252	0.689376	0.387181	0.118265
0.524016	0.539057	0.559501	0.424611
0.364240	0.707881	0.368965	0.345300
0.720254	0.518017	0.408374	0.238965
0.541362	0.606212	0.431139	0.330107
0.500451	0.584743	0.514882	0.313311
0.563683	0.711285	0.474227	0.465183
0.565374	0.497179	0.448769	0.300766
0.670367	0.649889	0.381539	0.437989
0.330120	0.598258	0.452806	0.217696
0.643262	0.423628	0.451488	0.429037
0.336383	0.638514	0.412625	0.269043
0.641518	0.557771	0.406588	0.523234
0.484462	0.297757	0.409613	0.406463
0.482366	0.526693	0.413265	0.423656
0.512033	0.669505	0.417390	0.197614
0.476083	0.508803	0.394663	0.357045
0.333372	0.302179	0.436092	0.370348
0.732748	0.508780	0.446511	0.610267
0.617068	0.452233	0.478107	0.382452
0.210447	0.470515	0.433979	0.250059
0.541835	0.373288	0.408689	0.415268
0.565113	0.348352	0.465581	0.463141
0.384680	0.451649	0.448793	0.140900
0.539277	0.769685	0.400437	0.408910
0.461752	0.463783	0.473103	0.303268
0.584231	0.517685	0.415986	0.249196
0.651084	0.804897	0.467982	0.512764
0.718360	0.631277	0.517953	0.588323
0.577288	0.590964	0.565910	0.347909
0.490538	0.484921	0.523945	0.472585
0.724895	0.361983	0.477862	0.500267
0.533684	0.490820	0.500375	0.315804
0.602166	0.463698	0.487679	0.430953
0.649157	0.348236	0.463698	0.515013
0.502681	0.497452	0.366456	0.390223
0.730910	0.524243	0.549617	0.385188
0.549681	0.402489	0.365369	0.498372
0.450400	0.352513	0.458557	0.345590
0.258640	0.325029	0.463237	0.276155
0.703291	0.493545	0.389676	0.310054
0.498359	0.561783	0.480819	0.381830
0.646611	0.692981	0.319708	0.234366
0.420435	0.506258	0.507634	0.409336
0.476490	0.299121	0.459066	0.433818
0.452731	0.342821	0.419262	0.341211
0.398222	0.460634	0.408163	0.317347
0.550729	0.475214	0.465883	0.342745
0.679130	0.684866	0.510998	0.558259
0.603142	0.685167	0.475636	0.473352
0.601056	0.413840	0.416911	0.331279
0.504125	0.500889	0.525777	0.088610
0.550544	0.450133	0.479004	0.474310
0.517735	0.559155	0.565170	0.377146
0.782382	0.318425	0.392880	0.643622
0.800777	0.682793	0.384140	0.452899
0.585186	0.254391	0.428368	0.457510
0.488395	0.644281	0.393751	0.332926
0.659319	0.502443	0.414258	0.417755
0.406677	0.574158	0.502014	0.174100
0.421331	0.410556	0.419997	0.410580
0.437801	0.562177	0.420230	0.343375
0.460973	0.539907	0.491469	0.407626
0.526147	0.412842	0.511513	0.290542
0.281033	0.382361	0.439431	0.285929
0.729311	0.516406	0.398324	0.615911
0.698815	0.618064	0.336403	0.332478
0.443594	0.527834	0.394687	0.412795
0.578929	0.425902	0.492812	0.536125
0.570700	0.787106	0.454262	0.307650
0.302791	0.644423	0.477921	0.279975
0.516532	0.584118	0.484369	0.314137
0.482108	0.425492	0.510989	0.481517
0.626346	0.363622	0.396756	0.560284
0.388157	0.309951	0.456285	0.299084
0.655970	0.496873	0.430317	0.427501
0.504534	0.337245	0.405284	0.415601
0.600438	0.445510	0.459712	0.339062
0.475068	0.439838	0.420736	0.423027
0.700297	0.617961	0.376302	0.342282
0.706666	0.748784	0.383854	0.255216
0.481655	0.530912	0.429565	0.456703
0.602443	0.618709	0.436614	0.510240
0.560667	0.586350	0.423774	0.494040
0.591716	0.437539	0.373471	0.227232
0.525405	0.382643	0.395954	0.503794
0.314749	0.667131	0.510884	0.236270
0.569562	0.451983	0.470359	0.262144
0.575612	0.689455	0.537018	0.431182
0.730600	0.506133	0.450421	0.457117
0.742627	0.627229	0.388579	0.432244
0.612088	0.457173	0.471319	0.394685
0.386482	0.756914	0.487885	0.344749
0.636763	0.529483	0.348473	0.517805
0.702465	0.461168	0.343809	0.500535
0.461061	0.517256	0.426028	0.448669
0.533878	0.463254	0.395887	0.428215
0.646699	0.514017	0.370990	0.331936
0.529226	0.588812	0.437292	0.429421
0.336913	0.593805	0.470150	0.202948
0.831752	0.537254	0.415048	0.339862
0.737556	0.685307	0.461912	0.359486
0.599394	0.777441	0.437147	0.416365
0.468448	0.494135	0.516281	0.291799
0.404949	0.586360	0.489240	0.216507
0.541416	0.497826	0.308759	0.344375
0.722527	0.515346	0.495502	0.611105
0.554173	0.457826	0.427382	0.346963
0.706954	0.449579	0.404962	0.532392
0.592945	0.453635	0.552566	0.407634
0.689785	0.477795	0.417704	0.361985
0.390920	0.565611	0.393946	0.384962
0.483215	0.693966	0.463359	0.409041
0.574009	0.460236	0.387657	0.508732
0.453547	0.449092	0.470886	0.332363
0.557164	0.524915	0.408533	0.295748
0.739660	0.747315	0.493997	0.264580
0.427138	0.709300	0.419573	0.291560
0.569806	0.568506	0.450273	0.370552
0.773461	0.377130	0.505871	0.423560
0.345929	0.477963	0.535342	0.362478
0.458678	0.556074	0.475725	0.102022
0.427263	0.389408	0.401364	0.438344
0.552151	0.414184	0.493942	0.438092
0.638856	0.634239	0.580617	0.342911
0.602853	0.573046	0.527378	0.515298
0.645017	0.536258	0.503929	0.161405
0.613280	0.608748	0.490896	0.203342
0.723413	0.441312	0.435720	0.487847
0.323551	0.454550	0.486720	0.338262
0.676145	0.550422	0.505041	0.424037
0.564187	0.549184	0.397614	0.414009
0.515746	0.504552	0.491859	0.405715
0.397746	0.425575	0.490960	0.256621
0.856661	0.509721	0.441774	0.550088
0.446074	0.582900	0.458142	0.317826
0.865936	0.549917	0.475934	0.496223
0.731406	0.514366	0.372238	0.528132
0.585521	0.590268	0.401306	0.460239
0.566411	0.497034	0.473449	0.445208
0.483410	0.476667	0.459473	0.256991
0.379490	0.218853	0.454863	0.336084
0.506421	0.532564	0.538786	0.322809
0.473273	0.613242	0.474573	0.397588
0.505334	0.573391	0.440258	0.471390
0.711272	0.454260	0.463133	0.516105
0.569113	0.483028	0.454433	0.277087
0.489124	0.783736	0.442474	0.298120
0.457113	0.455360	0.409123	0.354102
0.439847	0.408462	0.431317	0.315235
0.846648	0.593426	0.534653	0.281513
0.750205	0.485903	0.482119	0.624226
0.594622	0.473463	0.504244	0.431421
0.520297	0.682826	0.372701	0.425429
0.555526	0.431032	0.434578	0.209616
0.538872	0.586522	0.424105	0.380414
0.382311	0.396049	0.382777	0.293077
0.526732	0.673397	0.519025	0.429044
0.660906	0.528728	0.490746	0.448334
0.617510	0.447138	0.480378	0.502549
0.445021	0.692054	0.435579	0.230813
0.564262	0.528977	0.439477	0.441146
0.504446	0.375642	0.400598	0.397314
0.569411	0.403108	0.549187	0.484017
0.345460	0.694340	0.456509	0.333625
0.426556	0.477679	0.470037	0.295030
0.334587	0.417777	0.339847	0.379509
0.704221	0.385235	0.421565	0.362196
0.667433	0.355493	0.447221	0.435597
0.456060	0.623419	0.487452	0.407248
0.517474	0.337585	0.510336	0.317102
0.789580	0.503038	0.472653	0.397273
0.465358	0.609968	0.454950	0.422283
0.533239	0.630788	0.416792	0.245578
0.639323	0.578754	0.460931	0.429611
0.465337	0.385632	0.475145	0.289531
0.362155	0.638163	0.443897	0.325042
0.441269	0.369135	0.530620	0.344116
0.746018	0.475747	0.467543	0.398582
0.427954	0.550325	0.417464	0.424039
0.747822	0.525553	0.394403	0.259073
0.703495	0.645696	0.498842	0.505773
0.552370	0.654887	0.401883	0.259798
0.574111	0.488107	0.362418	0.272928
0.665087	0.457338	0.433865	0.415928
0.576354	0.463995	0.497821	0.477400
0.538087	0.582019	0.436161	0.375050
0.597624	0.609657	0.368716	0.396333
0.503158	0.319564	0.488113	0.403310
0.519571	0.417781	0.446219	0.406906
0.788840	0.243455	0.407668	0.417748
0.629184	0.501406	0.467151	0.445759
0.531545	0.505997	0.375970	0.292608
0.521246	0.524377	0.480125	0.387722
0.430497	0.400098	0.354851	0.421125
0.528237	0.504704	0.486765	0.449115
0.527361	0.512137	0.431045	0.483953
0.593366	0.232732	0.401132	0.491624
0.600140	0.457289	0.431535	0.518994
0.699135	0.445851	0.432816	0.433861
0.519878	0.530144	0.495638	0.451380
0.559971	0.654934	0.418569	0.432668
0.487106	0.553275	0.383692	0.265291
0.762047	0.517949	0.340026	0.499078
0.618557	0.669215	0.437055	0.332367
0.464652	0.463514	0.460038	0.440140
0.493404	0.550166	0.358154	0.442911
0.681329	0.687694	0.469409	0.544106
0.860198	0.470707	0.392514	0.593536
0.635927	0.301566	0.541162	0.439459
0.549941	0.592655	0.483322	0.472377
0.589599	0.368879	0.383967	0.421992
0.522768	0.561865	0.490169	0.482135
0.651470	0.548321	0.491607	0.560770
0.408450	0.621750	0.452139	0.291734
0.547633	0.726609	0.471733	0.363793
0.651016	0.692664	0.462762	0.445900
0.623234	0.760416	0.525863	0.315082
0.669107	0.280268	0.363523	0.589544
0.601241	0.624830	0.471375	0.384460
0.526652	0.707823	0.413786	0.427961
0.622986	0.262413	0.459685	0.564759
0.513743	0.523078	0.447251	0.190968
0.696144	0.667693	0.469759	0.471942
0.422286	0.575871	0.501148	0.358133
0.255571	0.584980	0.472778	0.300837
0.645747	0.513961	0.488988	0.439302
0.569870	0.516504	0.500568	0.436545
0.445536	0.604811	0.462375	0.223690
0.487978	0.611469	0.407961	0.246176
0.564330	0.610502	0.393259	0.450606
0.476595	0.485394	0.445529	0.384573
0.597057	0.521664	0.452652	0.370033
0.500876	0.533290	0.474913	0.373905
0.536863	0.657956	0.496553	0.304193
0.413563	0.569173	0.466234	0.358929
0.438813	0.437994	0.490027	0.441647
0.628830	0.412357	0.539887	0.563482
0.353910	0.266991	0.420653	0.402305
0.550457	0.490136	0.394358	0.508295
0.765963	0.646422	0.317767	0.381923
0.477413	0.410097	0.435923	0.375624
0.580899	0.324024	0.423589	0.545896
0.555579	0.647122	0.524374	0.416259
0.426888	0.424933	0.446837	0.117575
0.606349	0.548392	0.423519	0.292822
0.693295	0.363969	0.474549	0.243150
0.562989	0.417857	0.503749	0.504949
0.613943	0.597198	0.453621	0.393809
0.673562	0.428439	0.575342	0.434314
0.590438	0.367020	0.500965	0.460447
0.334396	0.604570	0.465084	0.333540
0.334719	0.533697	0.390632	0.331735
0.656628	0.428627	0.432592	0.531510
0.342943	0.623761	0.458740	0.342582
0.733962	0.602609	0.471461	0.569620
0.387211	0.401400	0.496478	0.358211
0.788581	0.352749	0.443607	0.611904
0.563853	0.514861	0.479829	0.214638
0.488343	0.512222	0.330727	0.451924
0.673297	0.792349	0.488814	0.413188
0.376134	0.568035	0.437354	0.231056
0.682009	0.465661	0.428304	0.513712
0.741026	0.521712	0.355606	0.318131
0.587373	0.556358	0.471495	0.496905
0.316589	0.534024	0.502941	0.264326
0.754766	0.570605	0.381362	0.364711
0.488039	0.531904	0.435913	0.438505
0.611361	0.543928	0.345589	0.430921
0.814479	0.457314	0.401562	0.445817
0.408519	0.391355	0.413096	0.341323
0.400697	0.462501	0.412403	0.290765
0.367294	0.563886	0.421868	0.379567
0.636560	0.544988	0.466302	0.516508
0.554365	0.518967	0.374977	0.262791
0.587780	0.333821	0.465369	0.452128
0.519085	0.523092	0.480266	0.430956
0.358288	0.574444	0.519468	0.240848
0.453992	0.503934	0.589590	0.274530
0.706423	0.546012	0.435860	0.554472
0.464659	0.514573	0.510083	0.352231
0.537768	0.355946	0.555442	0.418337
0.685650	0.671492	0.464303	0.561630
0.480007	0.414895	0.440165	0.462922
0.557424	0.712145	0.425230	0.353649
0.547828	0.479583	0.511965	0.259579
0.551291	0.559641	0.426195	0.456565
0.512718	0.593926	0.523933	0.395961
0.622994	0.462202	0.437565	0.372227
0.590766	0.528666	0.439208	0.358671
0.566579	0.529572	0.451511	0.339394
0.483171	0.312280	0.464718	0.383573
0.578241	0.516900	0.462156	0.346032
0.710190	0.525632	0.460285	0.535401
0.513050	0.549354	0.486642	0.374224
0.773146	0.572949	0.418350	0.582406
0.553409	0.342149	0.444260	0.470885
0.578644	0.479266	0.456302	0.401268
0.579452	0.637645	0.473258	0.423698
0.498353	0.488494	0.445182	0.337106
0.471915	0.544281	0.464509	0.335869
0.596472	0.600496	0.500779	0.363402
0.623745	0.486275	0.473569	0.425497
0.392447	0.321220	0.457220	0.324738
0.503317	0.600746	0.460886	0.369976
0.503823	0.540805	0.420099	0.365618
0.662004	0.576404	0.414674	0.511881
0.508692	0.530491	0.417428	0.330851
0.460761	0.283187	0.459560	0.346895
0.433481	0.626000	0.476689	0.398388
0.789459	0.785336	0.477313	0.391511
0.570575	0.670545	0.578766	0.355723
0.496245	0.317286	0.425034	0.326220
0.465528	0.630431	0.472085	0.381957
0.635382	0.854315	0.433484	0.367311
0.566292	0.683151	0.459429	0.310496
0.663887	0.578526	0.533956	0.383715
0.648592	0.695126	0.426866	0.501915
0.477482	0.585111	0.511666	0.306181
0.531581	0.540215	0.436471	0.423771
0.350353	0.417933	0.464308	0.397844
0.557060	0.567271	0.451787	0.432902
0.470861	0.524119	0.436656	0.421265
0.606239	0.463942	0.470697	0.517347
0.624177	0.338306	0.501169	0.578998
0.492411	0.510563	0.590779	0.420288
0.639091	0.363256	0.486211	0.424372
0.682611	0.348021	0.491841	0.435850
0.544771	0.704914	0.431883	0.470735
0.516877	0.529108	0.493873	0.472836
0.439911	0.454230	0.457208	0.264223
0.439555	0.387936	0.512698	0.450783
0.418274	0.289744	0.477346	0.407191
0.570249	0.480353	0.458304	0.520105
0.540872	0.478511	0.425607	0.386209
0.479943	0.789295	0.522013	0.382525
0.398132	0.491075	0.423915	0.396678
0.445677	0.312433	0.542390	0.411718
0.461869	0.474670	0.448874	0.245926
0.399269	0.540563	0.526676	0.344443
0.483943	0.375237	0.464372	0.451748
0.546933	0.507026	0.479848	0.274206
0.403028	0.545218	0.325475	0.197307
0.528428	0.560485	0.427193	0.350218
0.337838	0.371146	0.432283	0.273131
0.684808	0.443134	0.538523	0.386564
0.675439	0.721928	0.479246	0.541822
0.468772	0.725474	0.451340	0.391920
0.612830	0.744580	0.418357	0.470496
0.680670	0.473119	0.448510	0.422567
0.637815	0.546003	0.450892	0.424418
0.446825	0.493771	0.369352	0.447919
0.542345	0.515598	0.503857	0.401168
0.759569	0.607336	0.452159	0.363187
0.366804	0.470391	0.453679	0.400526
0.668569	0.590316	0.463935	0.484826
0.586924	0.387824	0.429794	0.351803
0.585501	0.719985	0.433733	0.442935
0.742983	0.534757	0.447590	0.535248
0.361096	0.654140	0.477834	0.344888
0.676783	0.439057	0.363752	0.399713
0.467781	0.425300	0.501794	0.422449
0.640274	0.609812	0.485872	0.354433
0.466508	0.471903	0.417834	0.441570
0.581391	0.544436	0.491112	0.312512
0.440680	0.414644	0.494793	0.433749
0.644419	0.791932	0.503303	0.375806
0.401843	0.469851	0.481306	0.312184
0.658051	0.343957	0.515340	0.433060
0.562447	0.505653	0.404748	0.338834
0.588832	0.568939	0.456144	0.393413
0.650081	0.580511	0.445170	0.297922
0.596612	0.594630	0.498590	0.489614
0.598590	0.401009	0.469135	0.416744
0.231137	0.533285	0.436170	0.289276
0.437962	0.707730	0.497974	0.364892
0.360079	0.585769	0.475208	0.304703
0.200705	0.619653	0.401302	0.279602
0.582283	0.618081	0.551328	0.477459
0.379637	0.808041	0.517493	0.281283
0.599285	0.477185	0.537908	0.443695
0.468181	0.669288	0.404774	0.371758
0.396385	0.475054	0.488539	0.306054
0.617901	0.719637	0.473567	0.411072
0.587235	0.355498	0.472069	0.523021
0.678841	0.675120	0.529249	0.385903
0.568401	0.599824	0.478536	0.272695
0.611620	0.341771	0.451691	0.217707
0.719826	0.635936	0.372608	0.575717
0.478013	0.616512	0.519499	0.363443
0.534995	0.490413	0.442236	0.273063
0.640113	0.576205	0.452432	0.434333
0.425234	0.532326	0.458242	0.420131
0.678405	0.356992	0.495008	0.446552
0.547557	0.288267	0.472398	0.519203
0.590210	0.614158	0.474479	0.437987
0.752288	0.378046	0.449576	0.503345
0.513870	0.541544	0.388119	0.344185
0.425867	0.386780	0.440465	0.453768
0.647944	0.614762	0.400748	0.431247
0.485441	0.528108	0.436779	0.411152
0.504364	0.453288	0.440236	0.333567
0.610891	0.628159	0.531991	0.485970
0.577666	0.703399	0.408216	0.447355
0.690881	0.592491	0.458042	0.470433
0.626080	0.728436	0.471444	0.489299
0.279718	0.483540	0.422767	0.329454
0.590532	0.460358	0.440767	0.469236
0.676678	0.759126	0.431147	0.528109
0.649317	0.518819	0.453856	0.301099
0.542179	0.601801	0.452086	0.227213
0.557796	0.657005	0.425802	0.424300
0.384513	0.374232	0.403987	0.145043
0.608497	0.650490	0.429039	0.435046
0.589115	0.685689	0.422641	0.160892
0.575997	0.557862	0.510699	0.512382
0.730741	0.289548	0.382188	0.440553
0.678815	0.627849	0.461784	0.361467
0.537837	0.437791	0.360349	0.246282
0.535828	0.347616	0.431282	0.397738
0.566779	0.465794	0.463759	0.395837
0.528734	0.244170	0.433750	0.398418
0.529943	0.463445	0.544067	0.482419
0.294806	0.433590	0.389011	0.319273
0.621866	0.586782	0.475041	0.485278
0.882388	0.477161	0.425349	0.649859
0.520277	0.666945	0.470459	0.233447
0.463364	0.532308	0.426034	0.443821
0.717970	0.462667	0.482634	0.314039
0.631625	0.435601	0.426930	0.504349
0.441103	0.360204	0.547763	0.354683
0.352792	0.592542	0.481123	0.278697
0.687702	0.417685	0.431380	0.411091
0.572463	0.423942	0.496860	0.490335
0.492767	0.378682	0.466881	0.349685
0.378125	0.471899	0.399683	0.374470
0.520051	0.580028	0.510087	0.330411
0.541811	0.381455	0.400646	0.268436
0.490949	0.661280	0.496130	0.176816
0.304735	0.391487	0.460684	0.379638
0.681149	0.399193	0.479614	0.430748
0.474371	0.805697	0.500354	0.301160
0.481129	0.571786	0.498494	0.453946
0.380714	0.484992	0.488917	0.367937
0.701389	0.402711	0.478111	0.543260
0.399045	0.614242	0.488731	0.398732
0.658013	0.528957	0.431171	0.255554
0.409780	0.342824	0.502438	0.386985
0.809584	0.407530	0.435648	0.570052
0.287661	0.401022	0.450703	0.369792
0.598300	0.437851	0.432935	0.331898
0.815344	0.427063	0.470324	0.553648
0.682188	0.683018	0.458636	0.416112
0.694111	0.620259	0.501050	0.418696
0.677819	0.550030	0.421754	0.479246
0.470453	0.503660	0.472283	0.384490
0.693224	0.654119	0.432752	0.506796
0.518557	0.251473	0.511318	0.468835
0.514858	0.365258	0.435108	0.250741
0.417425	0.568767	0.487243	0.293529
0.779643	0.574251	0.468333	0.485575
0.487497	0.581435	0.368224	0.321329
0.546821	0.280353	0.398606	0.483963
0.443081	0.429897	0.420701	0.420741
0.544868	0.587740	0.466527	0.481436
0.714450	0.762484	0.405561	0.469977
0.756158	0.615654	0.430096	0.508332
0.608545	0.443924	0.401962	0.489682
0.426333	0.479524	0.447205	0.428690
0.637893	0.246516	0.453979	0.479535
0.529813	0.513813	0.469150	0.446418
0.566018	0.392177	0.443216	0.465054
0.647536	0.382370	0.518464	0.481094
0.719829	0.571996	0.410040	0.222440
0.449912	0.696962	0.511516	0.291357
0.739782	0.694909	0.501564	0.467602
0.478400	0.515212	0.449670	0.318124
0.816569	0.457683	0.438000	0.578740
0.703650	0.470916	0.410404	0.383164
0.496389	0.391983	0.437775	0.482873
0.323014	0.625356	0.412205	0.306747
0.596017	0.555569	0.427654	0.387201
0.637554	0.440591	0.491048	0.515634
0.727333	0.253313	0.470695	0.389685
0.660690	0.467822	0.449784	0.436256
0.391490	0.523549	0.362783	0.369106
0.452568	0.543305	0.440420	0.331765
0.593581	0.652096	0.512088	0.462300
0.839225	0.594498	0.410151	0.094343
0.375702	0.476790	0.433063	0.392494
0.498339	0.487882	0.467149	0.383572
0.384321	0.466406	0.432724	0.281269
0.336173	0.553052	0.508827	0.312601
0.525703	0.480921	0.455057	0.469685
0.358969	0.227429	0.476257	0.379932
0.594405	0.319409	0.502152	0.279998
0.613637	0.517316	0.389094	0.385983
0.603917	0.559716	0.418941	0.368687
0.482398	0.375730	0.436437	0.466754
0.691720	0.157113	0.446303	0.264993
0.509654	0.463837	0.448657	0.306114
0.680081	0.412004	0.370697	0.541977
0.581766	0.261414	0.489014	0.460150
0.491884	0.501890	0.569058	0.425919
0.546462	0.514846	0.392271	0.401661
0.550278	0.375065	0.462808	0.462192
0.618306	0.436063	0.396308	0.451210
0.483594	0.424524	0.383605	0.399078
0.418531	0.400875	0.472140	0.297671
0.344246	0.505250	0.407889	0.309300
0.415639	0.440711	0.390926	0.356273
0.633410	0.639105	0.466475	0.479800
0.564228	0.294902	0.411818	0.304807
0.542870	0.530945	0.435261	0.477908
0.512800	0.710009	0.461583	0.392362
0.518911	0.601799	0.475360	0.466950
0.447424	0.520708	0.403807	0.365641
0.553624	0.584894	0.452333	0.453867
0.739957	0.399714	0.467014	0.296820
0.800281	0.353574	0.442932	0.557919
0.317914	0.516804	0.473897	0.326182
0.558840	0.606431	0.410502	0.426031
0.513540	0.521755	0.457870	0.443438
0.756854	0.342219	0.460464	0.619089
0.587730	0.499937	0.536567	0.101315
0.758188	0.539456	0.547076	0.396451
0.751641	0.622616	0.465176	0.557225
0.505847	0.460662	0.492215	0.325779
0.650791	0.447406	0.426433	0.434297
0.501410	0.423119	0.481067	0.457278
0.855606	0.584149	0.513770	0.529913
0.471240	0.603428	0.414395	0.265856
0.398360	0.555842	0.432147	0.406052
0.673035	0.407769	0.424826	0.404874
0.757608	0.243439	0.455748	0.497083
0.454741	0.579377	0.422447	0.207093
0.472966	0.644263	0.431523	0.312751
0.589928	0.486798	0.381366	0.425888
0.686968	0.593135	0.529939	0.503889
0.442619	0.679503	0.447743	0.206009
0.601382	0.320236	0.387855	0.448493
0.634618	0.562623	0.491301	0.541123
0.456673	0.349648	0.420319	0.473557
0.551803	0.659393	0.366156	0.294534
0.716968	0.739277	0.415932	0.427770
0.672400	0.476444	0.438469	0.427741
0.392304	0.317828	0.470354	0.409601
0.707052	0.608675	0.423158	0.580124
0.597732	0.359201	0.475580	0.301197
0.625334	0.526722	0.541150	0.505326
0.681554	0.515905	0.443873	0.345335
0.638312	0.565831	0.467127	0.455230
0.601202	0.557390	0.485896	0.340273
0.250839	0.291033	0.429756	0.224340
0.451787	0.539206	0.508886	0.141924
0.665881	0.432221	0.471973	0.559386
0.464848	0.563487	0.325067	0.182146
0.695143	0.345684	0.489181	0.563370
0.156027	0.393469	0.504177	0.237838
0.557315	0.322250	0.488481	0.450156
0.472986	0.435516	0.493343	0.367906
0.647046	0.537124	0.441198	0.466435
0.658149	0.501094	0.369897	0.209242
0.543886	0.656510	0.442921	0.468999
0.445425	0.897555	0.451707	0.341217
0.520505	0.523328	0.410210	0.434975
0.467610	0.509945	0.370561	0.414786
0.650798	0.635707	0.491459	0.424520
0.820922	0.358103	0.541686	0.567682
0.828964	0.395259	0.420764	0.233044
0.636117	0.480075	0.530391	0.459970
0.582454	0.230291	0.464278	0.532966
0.984896	0.601609	0.484738	0.513920
0.714781	0.555144	0.424137	0.578612
0.516194	0.493804	0.344249	0.414881
0.485602	0.620226	0.468044	0.345784
0.470190	0.471059	0.481333	0.409745
0.745626	0.533614	0.445238	0.395871
0.553669	0.562142	0.467469	0.471667
0.543083	0.682051	0.441100	0.440595
0.501387	0.620080	0.490999	0.322058
0.494752	0.516873	0.395273	0.453304
0.652998	0.449552	0.505623	0.443264
0.402119	0.375944	0.512198	0.422824
0.457901	0.457437	0.499742	0.149977
0.694920	0.507084	0.454793	0.380560
0.622101	0.569906	0.412695	0.508797
0.523713	0.445782	0.428346	0.406070
0.648132	0.740442	0.454254	0.438354
0.659604	0.464836	0.437201	0.357657
0.602276	0.498878	0.559294	0.198077
0.772097	0.416631	0.489908	0.477813
0.720677	0.633291	0.443093	0.307699
0.343981	0.608417	0.345737	0.309522
0.437433	0.353477	0.419620	0.377419
0.460781	0.359238	0.424508	0.437610
0.530356	0.606022	0.382150	0.463833
0.508324	0.653763	0.448300	0.442108
0.362756	0.352911	0.406502	0.329415
0.448572	0.303219	0.432095	0.413874
0.626345	0.305445	0.373233	0.525381
0.556696	0.398270	0.529825	0.344840
0.665544	0.311476	0.443344	0.416898
0.583049	0.259432	0.487852	0.362706
0.537666	0.405151	0.493106	0.250610
0.665476	0.417513	0.485899	0.382277
0.587228	0.548358	0.521616	0.380796
0.563624	0.552436	0.491916	0.460419
0.485251	0.361429	0.438962	0.475569
0.501925	0.527167	0.484274	0.392391
0.561343	0.644635	0.430238	0.453475
0.396740	0.612483	0.510018	0.376896
0.361610	0.473571	0.522999	0.267790
0.306228	0.357130	0.453750	0.258102
0.423366	0.742414	0.432514	0.371152
0.383463	0.414980	0.392025	0.302333
0.786195	0.616625	0.476317	0.396994
0.726657	0.577478	0.404238	0.550110
0.520398	0.419130	0.506481	0.311605
0.642055	0.274089	0.403781	0.434004
0.471124	0.375478	0.415399	0.269185
0.441670	0.726607	0.470815	0.355944
0.365388	0.631353	0.560650	0.353401
0.787462	0.449379	0.483025	0.522375
0.621490	0.355713	0.570863	0.549695
0.654817	0.717854	0.420766	0.373340
0.360288	0.450693	0.419904	0.381989
0.520957	0.603554	0.571822	0.332058
0.509015	0.289854	0.455980	0.504243
0.614904	0.453816	0.461328	0.258337
0.567782	0.230528	0.397443	0.402703
0.505672	0.536025	0.442351	0.327814
0.541539	0.363611	0.412897	0.483974
0.492222	0.274473	0.413161	0.457971
0.631635	0.555613	0.495790	0.310878
0.447608	0.387666	0.580549	0.176126
0.470637	0.382138	0.402882	0.370225
0.594342	0.380021	0.416486	0.444901
0.443596	0.421670	0.551106	0.331348
0.452907	0.815649	0.373066	0.395640
0.458746	0.352803	0.520068	0.356330
0.637691	0.674899	0.434275	0.532226
0.657812	0.621385	0.437711	0.520341
0.717191	0.443587	0.459323	0.621304
0.329321	0.539272	0.493120	0.156654
0.545385	0.506576	0.407930	0.296095
0.467180	0.691672	0.425335	0.415692
0.772391	0.626612	0.425718	0.403519
0.780935	0.410263	0.508978	0.517831
0.745313	0.625037	0.481675	0.493983
0.464058	0.615191	0.529751	0.292539
0.539408	0.355318	0.493457	0.411087
0.659885	0.456246	0.403461	0.450285
0.579126	0.527872	0.434925	0.354271
0.576737	0.446022	0.538927	0.178882
0.510633	0.482276	0.441146	0.422933
0.795372	0.430342	0.404163	0.531991
0.423750	0.266267	0.389271	0.438067
0.632093	0.504743	0.349563	0.511970
0.475809	0.500757	0.388088	0.323993
0.529891	0.571383	0.385063	0.340537
0.600387	0.874900	0.502475	0.432980
0.676066	0.426964	0.380397	0.585084
0.629535	0.579295	0.417971	0.444636
0.602781	0.489100	0.399046	0.295472
0.469293	0.405432	0.359936	0.293017
0.349258	0.354185	0.512826	0.161325
0.394053	0.469312	0.473740	0.205696
0.482523	0.545676	0.431155	0.457040
0.816879	0.431826	0.509151	0.661468
0.599770	0.449304	0.394448	0.444190
0.297835	0.567137	0.350593	0.266801
0.788447	0.598693	0.479003	0.340118
0.547668	0.460372	0.376500	0.481117
0.539303	0.622967	0.479314	0.091485
0.586732	0.764362	0.452142	0.431402
0.718740	0.673297	0.394459	0.449977
0.341229	0.538239	0.412946	0.247661
0.551837	0.371992	0.465826	0.429085
0.668583	0.711434	0.505056	0.350074
0.342445	0.457670	0.379869	0.391934
0.627816	0.466312	0.513618	0.387975
0.743941	0.464138	0.428542	0.316422
0.755027	0.585823	0.476817	0.375008
0.946057	0.494546	0.397185	0.647341
0.620565	0.402066	0.393034	0.291959
0.563331	0.346177	0.543225	0.272315
0.562042	0.722727	0.463022	0.364895
0.806873	0.435089	0.518614	0.613412
0.372202	0.680060	0.360863	0.302930
0.460395	0.665587	0.419362	0.419104
0.707822	0.415081	0.469989	0.587815
0.610490	0.670864	0.438170	0.337202
0.624880	0.435053	0.487546	0.321197
0.314841	0.673766	0.462738	0.322789
0.683099	0.279096	0.389140	0.312674
0.592356	0.713169	0.459604	0.325139
0.575694	0.513363	0.442256	0.323882
0.574689	0.583925	0.422057	0.482754
0.644033	0.621115	0.491871	0.452804
0.441276	0.420895	0.444959	0.437341
0.322192	0.488009	0.357754	0.211097
0.610584	0.606124	0.423257	0.485230
0.542912	0.387275	0.462629	0.477988
0.436389	0.499421	0.452080	0.430600
0.749961	0.760090	0.441054	0.438436
0.504124	0.385008	0.490432	0.384762
0.418549	0.526558	0.455517	0.269094
0.574978	0.715133	0.415168	0.335619
0.727407	0.751630	0.445864	0.489539
0.612900	0.478349	0.450958	0.404828
0.547942	0.486450	0.413703	0.499205
0.419809	0.609424	0.496018	0.381343
0.631567	0.611204	0.454868	0.531141
0.534534	0.191352	0.460743	0.517888
0.650856	0.306597	0.495895	0.405739
0.660388	0.510916	0.443580	0.500662
0.814973	0.552347	0.461334	0.376620
0.656345	0.638309	0.480499	0.418511
0.688185	0.565805	0.382990	0.466629
0.414278	0.567393	0.435559	0.413001
0.753917	0.500198	0.442066	0.562729
0.525577	0.413564	0.491707	0.307079
0.388621	0.663859	0.497011	0.218441
0.499488	0.494140	0.423708	0.435207
0.650664	0.565862	0.506709	0.456887
0.679898	0.553475	0.478092	0.402404
0.775827	0.652773	0.369633	0.190771
0.473524	0.541342	0.514068	0.388302
0.701625	0.545732	0.474124	0.318635
0.848759	0.624259	0.409701	0.492055
0.696295	0.503499	0.430456	0.496801
0.774018	0.468575	0.424462	0.295308
0.459667	0.437046	0.451622	0.456278
0.546329	0.640384	0.430873	0.368499
0.471219	0.276728	0.424270	0.479283
0.545143	0.669165	0.452561	0.285475
0.478384	0.526156	0.446998	0.378314
0.765456	0.504009	0.458263	0.423975
0.457637	0.494947	0.363473	0.409143
0.723967	0.717121	0.446560	0.530581
0.325593	0.511369	0.437223	0.305798
0.519933	0.591995	0.450832	0.311196
0.487818	0.481027	0.506716	0.282551
0.567358	0.505932	0.516197	0.369395
0.437763	0.575111	0.456546	0.219495
0.604774	0.669397	0.471581	0.443334
0.524299	0.635930	0.406385	0.454704
0.487029	0.558066	0.458161	0.452136
0.615873	0.440506	0.473947	0.469428
0.372955	0.236254	0.444795	0.416397
0.504790	0.521064	0.435232	0.307572
0.660194	0.472507	0.423405	0.514193
0.543577	0.319623	0.379806	0.536697
0.537925	0.540579	0.400292	0.479624
0.660695	0.544589	0.401730	0.469921
0.557189	0.575690	0.466649	0.360564
0.532680	0.398953	0.402879	0.227185
0.572480	0.275998	0.482334	0.428144
0.580889	0.244495	0.478284	0.463351
0.605257	0.553443	0.403452	0.339399
0.685008	0.731531	0.483100	0.469834
0.639723	0.614198	0.498272	0.535660
0.628539	0.634427	0.392400	0.464762
0.493829	0.582781	0.417126	0.356454
0.608479	0.672165	0.479522	0.395493
0.833940	0.597388	0.385613	0.464698
0.717614	0.532935	0.448080	0.582928
0.683175	0.626528	0.386309	0.392169
0.543763	0.472246	0.515703	0.374657
0.746315	0.136327	0.440244	0.549211
0.456757	0.461391	0.483900	0.391308
0.405193	0.548723	0.419791	0.334882
0.729840	0.552893	0.429902	0.269932
0.702573	0.678509	0.478218	0.495851
0.565101	0.679044	0.420469	0.461206
0.816258	0.175354	0.441215	0.644910
0.646898	0.766727	0.414470	0.474310
0.822011	0.533022	0.478953	0.541945
0.556924	0.493178	0.450707	0.358960
0.389103	0.457681	0.445823	0.218020
0.458182	0.628057	0.471531	0.272785
0.674254	0.511641	0.484193	0.314603
0.484283	0.360506	0.447931	0.374671
0.586523	0.576785	0.388950	0.254773
0.492063	0.514520	0.410790	0.348386
0.715253	0.559470	0.444974	0.440001
0.900251	0.705517	0.419539	0.212037
0.597248	0.613407	0.438360	0.384038
0.718891	0.461680	0.521703	0.442975
0.672682	0.605883	0.539341	0.526151
0.653008	0.349817	0.446774	0.382316
0.615171	0.554252	0.545156	0.409189
0.409850	0.411723	0.468193	0.351019
0.550112	0.413246	0.419389	0.452817
0.621588	0.718444	0.432985	0.425677
0.566420	0.392939	0.526725	0.297760
0.611386	0.477409	0.475234	0.417255
0.672059	0.544726	0.436235	0.378926
0.229444	0.504889	0.419488	0.314438
0.364205	0.547428	0.443746	0.286492
0.686503	0.735389	0.459465	0.338889
0.572841	0.274114	0.403353	0.365925
0.378886	0.585924	0.472129	0.381108
0.668655	0.605852	0.499178	0.556923
0.550876	0.401209	0.433069	0.415912
0.621230	0.602764	0.445807	0.463829
0.953714	0.631880	0.409632	0.313268
0.688887	0.751363	0.407696	0.350921
0.512355	0.563962	0.508740	0.371265
0.568734	0.483890	0.442547	0.398269
0.571814	0.471817	0.445233	0.229893
0.528956	0.397280	0.398549	0.132153
0.774074	0.449151	0.387581	0.606612
0.489720	0.702624	0.466514	0.361603
0.554621	0.560385	0.420867	0.307538
0.590778	0.435963	0.447599	0.150009
0.494112	0.397110	0.445581	0.492677
0.457678	0.594868	0.484303	0.246765
0.408442	0.494053	0.446278	0.417966
0.578929	0.501985	0.406026	0.356166
0.806641	0.567521	0.527529	0.348087
0.441897	0.705572	0.532530	0.334453
0.804695	0.706893	0.495400	0.358166
0.568043	0.239435	0.560377	0.225493
0.660692	0.545311	0.477932	0.395154
0.609053	0.471629	0.451785	0.326406
0.562225	0.506056	0.390732	0.468805
0.665228	0.414890	0.432670	0.425357
0.582708	0.767049	0.381414	0.341289
0.423903	0.425993	0.498279	0.258912
0.543798	0.672143	0.493654	0.427776
0.562054	0.399036	0.463249	0.441770
0.381655	0.502795	0.481397	0.366166
0.788674	0.503454	0.413298	0.391214
0.687551	0.686130	0.438314	0.346319
0.446794	0.544077	0.420128	0.378009
0.734581	0.643242	0.442687	0.489021
0.511505	0.642029	0.458219	0.453069
0.724320	0.431214	0.463401	0.364780
0.718624	0.488496	0.509816	0.437445
0.438659	0.587272	0.452155	0.412157
0.529670	0.384382	0.444161	0.422773
0.462187	0.471107	0.445424	0.238551
0.561414	0.679701	0.415669	0.382830
0.591414	0.528075	0.431432	0.484838
0.528264	0.558549	0.423690	0.365378
0.779566	0.325455	0.498777	0.416225
0.545716	0.346712	0.413339	0.501528
0.677689	0.462450	0.403788	0.333826
0.518755	0.684908	0.494743	0.407889
0.526157	0.494804	0.488161	0.473375
0.629232	0.503398	0.512135	0.448586
0.642954	0.439644	0.519554	0.369237
0.434450	0.284176	0.477041	0.472212
0.589471	0.452832	0.375872	0.383316
0.718815	0.620253	0.443926	0.567471
0.439748	0.573298	0.466560	0.371617
0.613362	0.696075	0.452862	0.412729
0.528761	0.586826	0.376574	0.418512
0.545684	0.704785	0.377338	0.374583
0.657989	0.519993	0.477950	0.344823
0.345650	0.483443	0.433402	0.353338
0.598769	0.475092	0.440779	0.474548
0.744475	0.563048	0.405669	0.426287
0.518522	0.319124	0.465427	0.233644
0.412776	0.468089	0.487648	0.417791
0.604530	0.640911	0.362325	0.311751
0.560452	0.671842	0.421692	0.264067
0.713297	0.261981	0.528418	0.416143
0.545255	0.819376	0.478689	0.334832
0.825292	0.554879	0.409793	0.394858
0.518305	0.369580	0.428349	0.502492
0.618094	0.593984	0.422572	0.331493
0.298427	0.676618	0.464906	0.264756
0.522900	0.721464	0.495131	0.405422
0.688348	0.437007	0.418816	0.384475
0.484941	0.472053	0.404719	0.448425
0.300617	0.433158	0.508654	0.362317
0.669395	0.424120	0.473554	0.544502
0.483257	0.522911	0.509905	0.371615
0.723240	0.396380	0.536407	0.606625
0.455898	0.413798	0.490403	0.434965
0.677183	0.406757	0.427328	0.539674
0.694848	0.679883	0.398223	0.454493
0.557578	0.502353	0.444802	0.436633
0.645341	0.472651	0.425083	0.236660
0.528058	0.723803	0.460374	0.368770
0.409892	0.417910	0.416895	0.435553
0.475828	0.550720	0.481452	0.390297
0.488941	0.548278	0.482387	0.458906
0.570398	0.615199	0.530463	0.451727
0.614164	0.387285	0.427206	0.563300
0.686157	0.421697	0.481932	0.376249
0.636206	0.558039	0.498172	0.380903
0.654853	0.518968	0.487061	0.490815
0.504753	0.630227	0.427799	0.287619
0.656698	0.347742	0.374770	0.391568
0.616727	0.507222	0.466528	0.489255
0.334979	0.649202	0.509451	0.349746
0.694893	0.485842	0.467901	0.523720
0.605784	0.731577	0.446803	0.398152
0.612487	0.695844	0.459224	0.489304
0.745394	0.396037	0.454798	0.490639
0.472079	0.635886	0.503366	0.339841
0.665837	0.584051	0.431011	0.369243
0.344803	0.459328	0.477384	0.209002
0.597626	0.570013	0.471781	0.425250
0.432564	0.633809	0.462787	0.335150
0.605658	0.509123	0.380507	0.422006
0.720579	0.300933	0.356183	0.386326
0.548837	0.511241	0.407586	0.437740
0.685726	0.650607	0.515358	0.505216
0.274376	0.313047	0.451548	0.346329
0.505479	0.315760	0.439812	0.438647
0.637477	0.622886	0.436035	0.368371
0.419569	0.509995	0.470968	0.311127
0.333528	0.582071	0.388656	0.267904
0.506482	0.635045	0.427614	0.455996
0.526015	0.489758	0.478979	0.444505
0.617874	0.519038	0.482098	0.336640
0.676995	0.477687	0.474225	0.449084
0.677872	0.456771	0.492377	0.561357
0.513419	0.645699	0.492214	0.452499
0.689074	0.670373	0.486897	0.432635
0.789614	0.625094	0.416215	0.473905
0.663744	0.532858	0.427639	0.340433
0.617687	0.653110	0.438686	0.402221
0.581167	0.661643	0.460814	0.467556
0.484956	0.338893	0.482698	0.395344
0.336556	0.525462	0.362613	0.330483
0.572732	0.659966	0.462007	0.320209
0.789458	0.380243	0.379839	0.307996
0.649838	0.440273	0.484563	0.474229
0.401954	0.509545	0.441146	0.219069
0.406827	0.548391	0.490379	0.383508
0.343250	0.412783	0.463745	0.337452
0.640490	0.514645	0.467795	0.271183
0.391743	0.654572	0.463067	0.140841
0.533557	0.593860	0.377153	0.142867
0.785985	0.604029	0.477568	0.457042
0.641330	0.468155	0.511542	0.496838
0.671435	0.653847	0.422078	0.453016
0.292112	0.563337	0.412234	0.344349
0.405299	0.593302	0.482847	0.305955
0.509182	0.485877	0.461313	0.476860
0.358060	0.418162	0.430274	0.355043
0.762443	0.417447	0.455581	0.464611
0.466282	0.555270	0.481548	0.307289
0.448629	0.565865	0.542426	0.319209
0.572261	0.500951	0.486919	0.475528
0.760403	0.627329	0.519382	0.496630
0.567674	0.600305	0.429147	0.250246
0.394768	0.448865	0.455888	0.386205
0.491265	0.735399	0.391932	0.304765
0.508114	0.506321	0.406858	0.476950
0.508890	0.453563	0.455176	0.411080
0.595122	0.432421	0.361178	0.368831
0.494788	0.419994	0.367027	0.317067
0.651086	0.567524	0.445698	0.486825
0.465200	0.352782	0.446530	0.374228
0.551582	0.451697	0.472515	0.467041
0.650984	0.738657	0.446328	0.428932
0.892653	0.535252	0.430492	0.287716
0.571276	0.522345	0.502764	0.501914
0.687293	0.563220	0.462006	0.548194
0.575152	0.679229	0.480938	0.348777
0.647875	0.574653	0.427346	0.402959
0.679820	0.656290	0.479735	0.545516
0.724446	0.590122	0.474945	0.287231
0.807455	0.521197	0.421388	0.342696
0.291787	0.537826	0.442534	0.208007
0.594655	0.486701	0.515585	0.461233
0.469749	0.376746	0.528712	0.126607
0.816078	0.640700	0.408253	0.469787
0.404437	0.506028	0.484550	0.377920
0.502197	0.458040	0.407137	0.358304
0.515082	0.327058	0.421604	0.444782
0.506565	0.451909	0.401412	0.336678
0.599910	0.361172	0.496829	0.414114
0.836279	0.302129	0.494655	0.335069
0.587279	0.417408	0.462084	0.407724
0.370069	0.467145	0.396368	0.395206
0.765836	0.502980	0.406743	0.496726
0.554329	0.592641	0.476157	0.329035
0.445628	0.215725	0.436057	0.379907
0.578495	0.669855	0.502668	0.210250
0.605371	0.536252	0.470868	0.271728
0.197543	0.449582	0.528944	0.194445
0.400615	0.529248	0.444295	0.278220
0.493901	0.782006	0.446818	0.413255
0.420338	0.550148	0.383188	0.316060
0.675926	0.418034	0.395224	0.581955
0.338952	0.611729	0.508524	0.360119
0.590686	0.638275	0.501647	0.317753
0.476922	0.529706	0.431733	0.265782
0.552824	0.628956	0.464074	0.381458
0.377918	0.340401	0.521724	0.430270
0.584673	0.562183	0.470001	0.211618
0.726836	0.598013	0.479100	0.439552
0.588099	0.372263	0.471157	0.335728
0.535484	0.382642	0.444038	0.424180
0.612426	0.458852	0.373359	0.413635
0.411869	0.416304	0.458353	0.422766
0.532324	0.331260	0.453237	0.265849
0.604925	0.625322	0.505432	0.508771
0.649375	0.681845	0.510253	0.346893
0.545735	0.528316	0.387700	0.482664
0.564735	0.543618	0.515876	0.431763
0.377024	0.420431	0.455422	0.306297
0.602767	0.524371	0.457707	0.495593
0.404257	0.608694	0.407563	0.386820
0.655049	0.417753	0.542589	0.541933
0.462663	0.379230	0.616271	0.374041
0.494489	0.861116	0.459613	0.385284
0.499299	0.478702	0.406638	0.411379
0.784282	0.579790	0.367388	0.485058
0.588766	0.611622	0.533521	0.497983
0.639200	0.455020	0.417113	0.460792
0.706398	0.654810	0.513044	0.444952
0.575858	0.509354	0.454836	0.476116
0.481751	0.665571	0.487117	0.275999
0.586107	0.462197	0.406315	0.314505
0.603738	0.523734	0.435296	0.266324
0.439146	0.552448	0.429746	0.147923
0.426868	0.550839	0.470925	0.240963
0.504347	0.528765	0.498314	0.396439
0.629022	0.331798	0.514130	0.279389
0.450968	0.621554	0.392731	0.368097
0.388940	0.547308	0.405288	0.358999
0.604233	0.464102	0.409163	0.496124
0.431850	0.554353	0.440019	0.333320
0.702659	0.268899	0.456827	0.215748
0.497388	0.471085	0.402452	0.432642
0.525042	0.640289	0.496081	0.196065
0.526428	0.522072	0.448999	0.464287
0.708048	0.589880	0.451139	0.504170
0.427603	0.441032	0.447575	0.402103
0.651429	0.466208	0.420221	0.357787
0.785724	0.585903	0.397513	0.365931
0.554774	0.517714	0.438659	0.507479
0.475698	0.611780	0.430028	0.260881
0.530321	0.641621	0.510893	0.461857
0.564335	0.492252	0.436083	0.454297
0.644213	0.695379	0.412622	0.524336
0.653207	0.606283	0.481788	0.361488
0.613586	0.379921	0.536367	0.486057
0.638901	0.437481	0.439068	0.341823
0.379790	0.367482	0.479020	0.317837
0.461484	0.349292	0.420382	0.460760
0.512297	0.311146	0.499119	0.479137
0.595037	0.565533	0.457452	0.507912
0.511251	0.444302	0.491488	0.493446
0.673843	0.531015	0.420648	0.437528
0.756310	0.595282	0.479321	0.439209
0.605913	0.361913	0.359253	0.551577
0.381182	0.320693	0.432315	0.266433
0.731930	0.455182	0.438171	0.512351
0.344653	0.593232	0.412587	0.297375
0.687477	0.384476	0.452304	0.310034
0.602832	0.688312	0.469798	0.403758
0.597896	0.593523	0.457878	0.363811
0.592891	0.589183	0.559099	0.499947
0.588761	0.553032	0.439204	0.245764
0.634128	0.386699	0.410610	0.284983
0.872299	0.436463	0.411432	0.383012
0.541454	0.536007	0.362850	0.195716
0.320244	0.328468	0.483793	0.343548
0.658251	0.561919	0.447139	0.276247
0.585627	0.614822	0.360203	0.290159
0.790392	0.518338	0.371950	0.164184
0.390123	0.843479	0.470897	0.318671
0.579534	0.479139	0.521267	0.420983
0.458560	0.529356	0.416774	0.286676
0.611635	0.670232	0.435521	0.514813
0.400889	0.663737	0.517003	0.365480
0.584367	0.550104	0.453105	0.474898
0.432937	0.452677	0.483610	0.425808
0.646720	0.242170	0.375997	0.602087
0.546731	0.396650	0.397622	0.424808
0.739430	0.316774	0.468653	0.356817
0.510114	0.669251	0.415773	0.446242
0.803131	0.379399	0.455912	0.492881
0.663466	0.260073	0.391442	0.469505
0.505722	0.467677	0.479177	0.482215
0.798342	0.438442	0.395900	0.562760
0.518064	0.706390	0.494822	0.381691
0.818151	0.355691	0.497609	0.582039
0.602400	0.425944	0.393302	0.376923
0.513685	0.423179	0.365114	0.360320
0.639530	0.465603	0.416772	0.382584
0.485055	0.656208	0.478503	0.359299
0.644247	0.692626	0.463837	0.341806
0.790877	0.668123	0.504967	0.425504
0.341676	0.585830	0.454021	0.336324
0.516845	0.633399	0.450691	0.450746
0.547019	0.482533	0.477979	0.410619
0.725312	0.417757	0.405505	0.599163
0.472707	0.222555	0.397479	0.427534
0.768493	0.510974	0.507994	0.595273
0.392378	0.430401	0.437487	0.299169
0.560244	0.649193	0.408189	0.382921
0.550604	0.548778	0.466374	0.385719
0.506455	0.754946	0.371414	0.339518
0.581929	0.409473	0.402639	0.532699
0.494397	0.584970	0.394990	0.344022
0.541298	0.406925	0.478036	0.460050
0.744550	0.555442	0.401112	0.515962
0.331290	0.565518	0.427783	0.307872
0.795537	0.461810	0.454786	0.411854
0.477039	0.286451	0.441345	0.171407
0.601927	0.423519	0.415599	0.552046
0.702756	0.441318	0.424742	0.481800
0.454832	0.579880	0.372831	0.355718
0.546185	0.676393	0.385119	0.326308
0.802995	0.586922	0.433132	0.531726
0.497771	0.493898	0.466712	0.457121
0.708648	0.385952	0.509943	0.563163
0.534268	0.448317	0.434776	0.167113
0.391321	0.366684	0.361181	0.368539
0.458692	0.454854	0.459650	0.453216
0.682802	0.750670	0.300783	0.408837
0.314891	0.439503	0.462519	0.318444
0.638148	0.574132	0.446235	0.497568
0.599893	0.491009	0.486986	0.296113
0.470473	0.610331	0.455572	0.323847
0.564657	0.507425	0.490602	0.398279
0.492559	0.372562	0.484614	0.238210
0.343025	0.476350	0.386571	0.326750
0.803169	0.442221	0.413293	0.551409
0.745289	0.460140	0.492274	0.521982
0.701967	0.536004	0.397635	0.585234
0.531078	0.681673	0.488860	0.328236
0.584670	0.639595	0.425693	0.399399
0.306361	0.737921	0.365176	0.292351
0.763986	0.323482	0.460537	0.535717
0.741682	0.501056	0.469141	0.408579
0.579070	0.614730	0.405958	0.479560
0.524220	0.506949	0.447364	0.344749
0.427215	0.457451	0.435646	0.439394
0.843404	0.593296	0.436939	0.634731
0.441872	0.418933	0.539074	0.442692
0.493116	0.598143	0.504182	0.384101
0.692549	0.498836	0.514174	0.520781
0.540646	0.537492	0.442422	0.316442
0.741676	0.540785	0.476130	0.597144
0.683112	0.381497	0.388599	0.337197
0.275729	0.315282	0.507471	0.167146
0.663086	0.677017	0.453561	0.388077
0.536762	0.543738	0.549909	0.387884
0.653163	0.474877	0.375592	0.379680
0.716040	0.380376	0.409305	0.561275
0.275896	0.380256	0.498712	0.239640
0.413079	0.392880	0.605528	0.430135
0.543875	0.644836	0.455980	0.345248
0.378435	0.640283	0.399726	0.252808
0.429287	0.609562	0.479129	0.414220
0.630963	0.593038	0.424867	0.353980
0.621260	0.634034	0.484346	0.458281
0.716453	0.610687	0.468113	0.390443
0.553482	0.767068	0.412999	0.374270
0.455044	0.525496	0.487667	0.395082
0.424604	0.000000	0.435589	0.446127
0.804503	0.585203	0.466341	0.399306
0.264521	0.504052	0.499403	0.337512
0.586546	0.599509	0.510320	0.241954
0.305498	0.443013	0.425457	0.343413
0.584242	0.560311	0.452824	0.405553
0.638618	0.491963	0.535863	0.234084
0.519037	0.561474	0.428288	0.396723
0.541208	0.335115	0.410480	0.382765
0.762093	0.732834	0.437761	0.454369
0.348218	0.448394	0.379924	0.366124
0.575244	0.366362	0.473648	0.379727
0.660149	0.534667	0.463723	0.394558
0.561637	0.577786	0.467766	0.486188
0.453388	0.393469	0.478233	0.426964
0.138639	0.576440	0.502590	0.224255
0.353376	0.692987	0.465154	0.304670
0.776903	0.702390	0.414727	0.433806
0.672851	0.495691	0.390870	0.477772
0.527869	0.383526	0.450283	0.339581
0.733360	0.379701	0.468196	0.628553
0.645135	0.508147	0.411103	0.402635
0.578008	0.843997	0.347840	0.437435
0.569362	0.399017	0.380096	0.476549
0.805173	0.684604	0.445910	0.456622
0.685057	0.558292	0.445384	0.420753
0.485909	0.426956	0.448853	0.363651
0.487928	0.490281	0.518911	0.418735
0.292858	0.465865	0.509068	0.235673
0.416985	0.665274	0.362550	0.392597
0.549664	0.512364	0.414028	0.406553
0.676877	0.601407	0.458777	0.425999
0.489468	0.261730	0.469130	0.351513
0.304736	0.578546	0.460956	0.189939
0.450269	0.612206	0.440120	0.424495
0.259851	0.554166	0.410015	0.314648
0.574253	0.647189	0.416382	0.356835
0.761411	0.560937	0.473215	0.531989
0.517810	0.600444	0.425663	0.441354
0.432688	0.399456	0.469542	0.284840
0.251818	0.418756	0.437712	0.324111
0.594971	0.484147	0.415288	0.328385
0.560867	0.484779	0.429133	0.257287
0.553810	0.521323	0.454483	0.276094
0.715196	0.659889	0.435585	0.301662
0.431752	0.461737	0.500174	0.443398
0.743822	0.477222	0.489551	0.463364
0.566863	0.542425	0.466822	0.370283
0.465250	0.467146	0.445880	0.439857
0.599504	0.624543	0.425898	0.328892
0.481963	0.351991	0.385267	0.430973
0.467506	0.458654	0.395545	0.338477
0.529449	0.347766	0.404150	0.441316
0.501956	0.625760	0.411531	0.384358
0.563599	0.647950	0.454910	0.466725
0.343719	0.315286	0.469617	0.324258
0.641384	0.707028	0.422389	0.484070
0.308544	0.652666	0.525988	0.298357
0.602157	0.604264	0.462315	0.442803
0.774039	0.545874	0.399033	0.560953
0.601737	0.461879	0.431098	0.429843
0.405083	0.438336	0.500934	0.375460
0.481983	0.356140	0.388301	0.441645
0.565181	0.455055	0.455665	0.517298
0.451450	0.687806	0.441160	0.278044
0.469157	0.461405	0.441930	0.465185
0.258844	0.581555	0.543005	0.317909
0.460254	0.591664	0.427733	0.441247
0.591013	0.312776	0.422033	0.431930
0.801671	0.602542	0.513290	0.420170
0.595192	0.584501	0.442273	0.466410
0.715824	0.411817	0.465978	0.509512
0.358140	0.588276	0.379507	0.143800
0.573516	0.353150	0.456790	0.406330
0.245415	0.643801	0.494867	0.000000
0.446368	0.338224	0.465153	0.401555
0.645564	0.550502	0.350798	0.403994
0.728431	0.486601	0.416921	0.544255
0.259500	0.489839	0.489510	0.306027
0.405689	0.638816	0.477969	0.324571
0.842673	0.612763	0.493613	0.381531
0.728424	0.531102	0.495171	0.511356
0.604058	0.645924	0.447747	0.342091
0.771489	0.485809	0.341303	0.543727
0.707886	0.553697	0.588128	0.451521
0.385066	0.483660	0.424826	0.323012
0.512086	0.820530	0.425694	0.403496
0.527269	0.480777	0.441641	0.380911
0.474853	0.423044	0.451964	0.382082
0.517528	0.513600	0.478629	0.419020
0.514430	0.487389	0.500595	0.296030
0.602889	0.420417	0.526120	0.377514
0.520353	0.483510	0.499071	0.420263
0.785690	0.584724	0.499540	0.554467
0.661249	0.582548	0.458784	0.490892
0.615196	0.720325	0.438681	0.393103
0.691394	0.543244	0.406682	0.363579
0.564287	0.539561	0.457551	0.349005
0.835136	0.476163	0.483499	0.410255
0.499851	0.482929	0.485467	0.284037
0.634731	0.518667	0.404536	0.465226
0.688152	0.846681	0.419949	0.302281
0.530362	0.489835	0.500122	0.311948
0.734322	0.447926	0.475338	0.386261
0.499881	0.577307	0.509019	0.423436
0.546850	0.411067	0.548292	0.518940
0.461829	0.383584	0.410818	0.343832
0.405633	0.563795	0.342523	0.126103
0.853077	0.549974	0.433841	0.518905
0.535129	0.314384	0.438522	0.364825
0.669081	0.544148	0.460564	0.299275
0.412817	0.483039	0.506781	0.320082
0.491401	0.514487	0.471119	0.213919
0.550446	0.482283	0.460485	0.452764
0.643039	0.563665	0.440918	0.367720
0.750631	0.633804	0.446344	0.549351
0.727434	0.576432	0.413292	0.310481
0.533351	0.722243	0.402861	0.441272
0.198500	0.445860	0.416722	0.283489
0.609266	0.445942	0.448467	0.307674
0.476357	0.449012	0.474581	0.432649
0.556923	0.699315	0.442809	0.470874
0.592308	0.408160	0.551459	0.502784
0.342098	0.397735	0.420052	0.285232
0.589890	0.561650	0.446325	0.504917
0.559138	0.432330	0.488213	0.492670
0.763378	0.527807	0.429374	0.305346
0.637856	0.490701	0.485805	0.516246
0.575205	0.587968	0.412746	0.449533
0.386151	0.317429	0.462313	0.439713
0.342984	0.490120	0.443734	0.268113
0.518185	0.502077	0.443035	0.250437
0.415807	0.684018	0.546128	0.375175
0.487596	0.639974	0.411880	0.443916
0.509810	0.517431	0.494158	0.454512
0.534036	0.434300	0.434479	0.384292
0.609681	0.320167	0.513051	0.451919
0.557176	0.556989	0.366794	0.390906
0.401340	0.537771	0.437940	0.383158
0.592284	0.423178	0.510499	0.362622
0.638792	0.449532	0.424822	0.498543
0.441765	0.583982	0.414516	0.414202
0.511884	0.314699	0.325412	0.446115
0.494402	0.546813	0.412590	0.454053
0.788463	0.464207	0.465404	0.327359
0.749561	0.483331	0.428038	0.207501
0.569501	0.513204	0.434032	0.251877
0.605993	0.366659	0.383604	0.430150
0.412068	0.633647	0.470204	0.183382
0.437525	0.479287	0.467242	0.410004
0.602746	0.396035	0.455315	0.401956
0.657578	0.502026	0.444184	0.263332
0.468439	0.567070	0.471130	0.333536
0.363394	0.372087	0.412236	0.385781
0.443130	0.477517	0.449187	0.425758
0.217710	0.445588	0.413006	0.318684
0.551225	0.391146	0.478265	0.483939
0.630369	0.520857	0.513654	0.238891
0.719942	0.429319	0.467367	0.520993
0.539636	0.399756	0.435750	0.419403
0.759182	0.548371	0.475967	0.383385
0.617244	0.661884	0.422011	0.500980
0.607837	0.554246	0.476795	0.405717
0.352368	0.482171	0.424542	0.358485
0.446293	0.465271	0.489118	0.454270
0.720520	0.291123	0.451022	0.629901
0.520192	0.590559	0.519578	0.283458
0.671501	0.403245	0.471468	0.597620
0.480412	0.255042	0.564205	0.426347
0.598586	0.635714	0.502982	0.430948
0.482280	0.522981	0.371414	0.459830
0.733239	0.526706	0.432381	0.442310
0.574073	0.675150	0.430344	0.125064
0.671408	0.456842	0.537959	0.409481
0.571957	0.620444	0.417434	0.341464
0.425581	0.347228	0.438426	0.327831
0.381074	0.459418	0.436230	0.376397
0.733321	0.619473	0.507338	0.311266
0.439553	0.331328	0.463680	0.464829
0.589215	0.315040	0.380173	0.499727
0.644974	0.412149	0.424259	0.455280
0.601053	0.658767	0.416464	0.352585
0.724536	0.597283	0.386638	0.471482
0.652598	0.363367	0.445823	0.343660
0.484149	0.633974	0.499268	0.441920
0.678959	0.423441	0.498181	0.575044
0.694384	0.397143	0.485792	0.567189
0.613488	0.687337	0.366498	0.405041
0.390942	0.189254	0.411695	0.310626
0.478899	0.593958	0.434974	0.254291
0.699199	0.468449	0.479408	0.509534
0.514372	0.709586	0.424011	0.364011
0.303764	0.518680	0.529099	0.295469
0.509271	0.418647	0.299760	0.383197
0.687136	0.624770	0.444766	0.346786
0.576694	0.558310	0.475714	0.484883
0.493664	0.637406	0.355296	0.418531
0.553847	0.604609	0.414430	0.477968
0.497913	0.597499	0.342090	0.409498
0.593814	0.359457	0.477249	0.535535
0.622466	0.512819	0.392315	0.430826
0.686927	0.500501	0.421931	0.499063
0.299863	0.451900	0.454403	0.304670
0.383398	0.425124	0.488478	0.311830
0.659882	0.599621	0.463416	0.454385
0.694938	0.371563	0.423878	0.244413
0.600928	0.425794	0.391550	0.351080
0.722272	0.561867	0.413349	0.210992
0.633041	0.560926	0.463879	0.320023
0.676330	0.451335	0.546246	0.495026
0.390886	0.566182	0.527409	0.355196
0.423767	0.706507	0.471056	0.374312
0.354969	0.448908	0.459664	0.401315
0.549858	0.583897	0.388179	0.385138
0.579188	0.592562	0.412744	0.490882
0.712661	0.675588	0.403480	0.220657
0.608969	0.511204	0.420165	0.375198
0.439371	0.494488	0.448515	0.445062
0.450233	0.377400	0.381025	0.302607
0.522434	0.604500	0.378453	0.467035
0.544648	0.245149	0.458734	0.415015
0.403805	0.583011	0.411921	0.361771
0.414555	0.316387	0.426370	0.393796
0.512223	0.507705	0.456338	0.376224
0.380508	0.598413	0.403178	0.234631
0.550804	0.486171	0.467213	0.509407
0.582959	0.363521	0.417354	0.406314
0.473328	0.534127	0.445964	0.427076
0.665487	0.493661	0.515912	0.580059
0.429720	0.573796	0.478070	0.323278
0.719890	0.621447	0.478691	0.385142
0.605445	0.502898	0.383521	0.376695
0.350382	0.398060	0.396621	0.399273
0.673913	0.468115	0.420329	0.273091
0.725016	0.422586	0.544575	0.263958
0.452740	0.545757	0.421963	0.379982
0.677222	0.568083	0.465924	0.558220
0.666542	0.598460	0.428965	0.420137
0.503876	0.514333	0.430630	0.348698
0.531221	0.570731	0.504075	0.309345
0.539240	0.404937	0.501660	0.513808
0.449674	0.591794	0.499515	0.287324
0.297375	0.627702	0.436318	0.276526
0.658568	0.584773	0.384474	0.515295
0.525019	0.782262	0.478924	0.290399
0.733509	0.693666	0.399635	0.388818
0.691801	0.534616	0.450517	0.486400
0.835021	0.434833	0.463707	0.569810
0.739882	0.624828	0.456293	0.495267
0.530365	0.412154	0.381546	0.345057
0.571915	0.550464	0.557911	0.479210
0.502569	0.419593	0.542378	0.412009
0.577658	0.590067	0.494367	0.343905
0.507848	0.338404	0.371927	0.401296
0.603846	0.203797	0.450846	0.563522
0.422000	0.369876	0.473462	0.455372
0.754825	0.356711	0.475249	0.418595
0.466058	0.527905	0.443254	0.442707
0.309632	0.603576	0.453613	0.233884
0.797115	0.537651	0.475806	0.577985
0.573564	0.519448	0.506436	0.198743
0.563493	0.650446	0.412795	0.274554
0.697415	0.377969	0.423755	0.532781
0.590855	0.436064	0.437238	0.376533
0.611298	0.470728	0.345360	0.442787
0.548506	0.567791	0.513746	0.449817
0.321604	0.676492	0.467671	0.318557
0.374152	0.442757	0.446369	0.326104
0.457702	0.672349	0.534468	0.425386
0.508701	0.415712	0.473492	0.491150
0.474555	0.235180	0.442188	0.383276
0.530266	0.418119	0.375900	0.423441
0.525111	0.515923	0.434393	0.481328
0.718326	0.629791	0.494020	0.374999
0.507877	0.638556	0.475605	0.434780
0.418386	0.402307	0.349129	0.370622
0.401207	0.347944	0.417320	0.290770
0.416813	0.563055	0.396863	0.289594
0.623623	0.490714	0.524768	0.442543
0.771486	0.571681	0.408020	0.243491
0.545593	0.624385	0.526618	0.465961
0.738403	0.340862	0.516692	0.366948
0.374718	0.486501	0.477476	0.335731
0.491176	0.431665	0.391181	0.358921
0.352830	0.570017	0.422955	0.357289
0.486460	0.343946	0.418370	0.382677
0.691292	0.712944	0.492294	0.446727
0.570583	0.499884	0.389046	0.463893
0.411486	0.425541	0.468917	0.400649
0.353782	0.312636	0.442330	0.250786
0.698307	0.454664	0.490605	0.416859
0.430501	0.436750	0.525978	0.298205
0.711284	0.444371	0.404751	0.370656
0.314569	0.436011	0.529065	0.323515
0.349778	0.460101	0.398721	0.265004
0.727946	0.490046	0.502792	0.447996
0.481660	0.673535	0.481451	0.367814
0.755534	0.622301	0.379869	0.446803
0.303153	0.428759	0.470012	0.366360
0.735631	0.316732	0.445812	0.509293
0.736954	0.762903	0.388240	0.434037
0.588545	0.648683	0.422159	0.344665
0.519314	0.313904	0.368669	0.454002
0.555371	0.356232	0.383286	0.467017
0.571991	0.402193	0.434859	0.465862
0.605544	0.478621	0.430562	0.476588
0.341758	0.568661	0.454818	0.323662
0.365589	0.342238	0.384059	0.400952
0.482371	0.282452	0.413719	0.255657
0.476801	0.333119	0.449342	0.464443
0.682320	0.603024	0.467403	0.396477
0.621200	0.662610	0.392922	0.512203
0.565341	0.632290	0.492160	0.419987
0.384062	0.604812	0.425491	0.214999
0.601786	0.590120	0.416547	0.524546
0.283200	0.716146	0.474689	0.219273
0.663759	0.581892	0.510010	0.529536
0.521230	0.670622	0.380815	0.347716
0.520581	0.314747	0.440456	0.420760
0.612600	0.597380	0.436412	0.460828
0.555888	0.663622	0.463755	0.483222
0.638973	0.408963	0.405957	0.378897
0.504791	0.695171	0.432859	0.438587
0.536817	0.540818	0.453661	0.450872
0.705450	0.485495	0.500769	0.276766
0.721110	0.673702	0.424843	0.447228
0.628218	0.561911	0.460489	0.496501
0.413824	0.314821	0.457012	0.395076
0.443424	0.623257	0.491591	0.333184
0.491825	0.453934	0.413127	0.442420
0.627068	0.722978	0.515734	0.346151
0.538676	0.630902	0.456877	0.470511
0.738116	0.623470	0.454965	0.156401
0.655388	0.567086	0.440347	0.327497
0.371712	0.336835	0.435446	0.365863
0.624985	0.641480	0.520412	0.458195
0.413512	0.672900	0.381250	0.265382
0.810095	0.666545	0.389098	0.474822
0.643710	0.411970	0.373467	0.405389
0.609784	0.464012	0.463604	0.512813
0.745051	0.557487	0.483274	0.441680
0.644871	0.594386	0.477486	0.433918
0.538586	0.521069	0.404034	0.389800
0.563732	0.551927	0.420787	0.417718
0.629038	0.385050	0.454642	0.305839
0.630276	0.550121	0.326023	0.421304
0.463373	0.257897	0.359168	0.490798
0.555392	0.660232	0.412447	0.432286
0.630355	0.599230	0.492998	0.394185
0.617196	0.604164	0.426060	0.341530
0.545598	0.460056	0.433671	0.477992
0.728016	0.646193	0.471938	0.479047
0.463271	0.474587	0.491928	0.266511
0.566938	0.408353	0.525320	0.207441
0.655475	0.634409	0.479483	0.475902
0.531077	0.479250	0.433616	0.314433
0.427210	0.622348	0.496324	0.313011
0.551118	0.531313	0.475379	0.324086
0.406815	0.374717	0.461485	0.200849
0.578269	0.476723	0.484639	0.482688
0.283416	0.450817	0.424257	0.356350
0.565202	0.658755	0.403216	0.117543
0.642951	0.562491	0.463134	0.401287
0.345305	0.536728	0.449932	0.316704
0.518956	0.251926	0.438955	0.419461
0.511449	0.379715	0.450910	0.456293
0.715802	0.347264	0.417241	0.390983
0.225338	0.344557	0.406234	0.332879
0.535004	0.423687	0.449960	0.464221
0.572037	0.411368	0.505750	0.537149
0.408988	0.816077	0.432940	0.331102
0.580636	0.395304	0.459432	0.530637
0.617668	0.467541	0.457266	0.544157
0.599785	0.553896	0.411260	0.300545
0.768024	0.500996	0.469621	0.307983
0.510298	0.731802	0.344816	0.372418
0.494117	0.515462	0.453692	0.469268
0.499109	0.837900	0.457381	0.374987
0.478231	0.402595	0.450037	0.474637
0.421641	0.609186	0.411430	0.400166
0.751180	0.518921	0.515898	0.397263
0.611021	0.377148	0.500028	0.468496
0.777458	0.254763	0.367163	0.516631
0.530072	0.395971	0.464462	0.480268
0.502407	0.582008	0.465888	0.399658
0.494431	0.428195	0.512007	0.415226
0.344451	0.616737	0.510599	0.233596
0.575013	0.757433	0.439421	0.377350
0.555695	0.567894	0.454934	0.422903
0.692375	0.476992	0.451450	0.494920
0.600295	0.429698	0.530800	0.518039
0.607495	0.435114	0.442345	0.370556
0.516618	0.542270	0.488240	0.352892
0.296600	0.391704	0.460731	0.311558
0.354521	0.436370	0.448551	0.399703
0.608524	0.428974	0.385369	0.313728
0.594927	0.593286	0.537531	0.316182
0.626189	0.531345	0.456228	0.516205
0.512978	0.405549	0.427813	0.497801
0.650483	0.622109	0.468259	0.479881
0.297613	0.560955	0.463595	0.275354
0.454449	0.407703	0.400135	0.424524
0.603790	0.679077	0.449629	0.401731
0.621818	0.580760	0.470967	0.352532
0.415895	0.438620	0.451586	0.288714
0.713682	0.687595	0.446464	0.275831
0.511568	0.450926	0.392278	0.371849
0.640619	0.356621	0.455612	0.470523
0.437001	0.525012	0.440757	0.376335
0.476676	0.477979	0.446410	0.419964
0.827576	0.608171	0.457760	0.561605
0.567755	0.611218	0.440303	0.368996
0.513648	0.482209	0.473997	0.372958
0.603663	0.456925	0.505755	0.369628
0.674703	0.394167	0.386982	0.510563
0.491575	0.368473	0.404875	0.492126
0.595735	0.675334	0.510434	0.349628
0.546015	0.624694	0.532651	0.433781
0.647886	0.247958	0.376663	0.461565
0.609428	0.394855	0.456263	0.439809
0.718190	0.832339	0.426296	0.400376
0.462535	0.514574	0.440444	0.443260
0.584825	0.582765	0.469501	0.375336
0.612932	0.581529	0.516944	0.458711
0.358022	0.742460	0.410546	0.207091
0.612924	0.637133	0.489214	0.417351
0.381237	0.578566	0.423096	0.390558
0.487583	0.525445	0.451600	0.285070
0.836195	0.342420	0.484557	0.669913
0.415034	0.240991	0.386095	0.422502
0.573219	0.498263	0.475432	0.342574
0.829652	0.685285	0.429105	0.308954
0.871622	0.414488	0.566413	0.591732
0.604913	0.571712	0.458887	0.299547
0.462240	0.446447	0.401614	0.346960
0.491868	0.551731	0.381295	0.353614
0.606339	0.507673	0.462456	0.254064
0.455011	0.594066	0.395648	0.437550
0.409560	0.681896	0.472563	0.382231
0.432954	0.721426	0.413830	0.337527
0.918714	0.473553	0.437354	0.513931
0.303073	0.426200	0.504258	0.332157
0.406521	0.551273	0.456909	0.368559
0.516483	0.474602	0.491242	0.417263
0.799299	0.421638	0.505437	0.349957
0.715586	0.341250	0.463068	0.534177
0.374889	0.320222	0.471322	0.305580
0.736510	0.456885	0.439319	0.483800
0.548275	0.647146	0.436559	0.373917
0.599194	0.717731	0.340637	0.387697
0.626518	0.416266	0.406399	0.529148
0.400317	0.426610	0.414969	0.362639
0.429848	0.414845	0.451816	0.451061
0.818455	0.417961	0.416652	0.381466
0.644069	0.559050	0.468961	0.282506
0.607952	0.681479	0.492133	0.304129
0.870937	0.358448	0.407895	0.325533
0.692505	0.649422	0.403923	0.462492
0.657887	0.527809	0.426607	0.440432
0.304255	0.515437	0.458319	0.286597
0.375971	0.487290	0.453502	0.357901
0.536101	0.457090	0.466648	0.399280
0.602318	0.561200	0.505042	0.485248
0.747561	0.638005	0.409368	0.394089
0.462150	0.479115	0.433226	0.278074
0.499386	0.261686	0.476471	0.510306
0.466389	0.508703	0.479109	0.328591
0.445933	0.552331	0.454301	0.207973
0.553755	0.607423	0.407868	0.308118
0.634500	0.459887	0.411737	0.391031
